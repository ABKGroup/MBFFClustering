VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_160x118
  FOREIGN fakeram7_160x118 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 15.390 BY 42.000 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.192 0.024 0.216 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.288 0.024 0.312 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.384 0.024 0.408 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.480 0.024 0.504 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.576 0.024 0.600 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.672 0.024 0.696 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.768 0.024 0.792 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.864 0.024 0.888 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.960 0.024 0.984 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.056 0.024 1.080 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.152 0.024 1.176 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.344 0.024 1.368 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.536 0.024 1.560 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.632 0.024 1.656 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.728 0.024 1.752 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.920 0.024 1.944 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.016 0.024 2.040 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.112 0.024 2.136 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.208 0.024 2.232 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.304 0.024 2.328 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.400 0.024 2.424 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.496 0.024 2.520 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.592 0.024 2.616 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.688 0.024 2.712 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.784 0.024 2.808 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.880 0.024 2.904 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.976 0.024 3.000 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.072 0.024 3.096 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.264 0.024 3.288 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.360 0.024 3.384 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.456 0.024 3.480 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.552 0.024 3.576 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.648 0.024 3.672 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.744 0.024 3.768 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.840 0.024 3.864 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.936 0.024 3.960 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.032 0.024 4.056 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.224 0.024 4.248 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.320 0.024 4.344 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.416 0.024 4.440 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.512 0.024 4.536 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.608 0.024 4.632 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.704 0.024 4.728 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.800 0.024 4.824 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.992 0.024 5.016 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.088 0.024 5.112 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.184 0.024 5.208 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.280 0.024 5.304 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.376 0.024 5.400 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.568 0.024 5.592 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.664 0.024 5.688 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.760 0.024 5.784 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.856 0.024 5.880 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.952 0.024 5.976 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 0.024 6.072 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.144 0.024 6.168 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.240 0.024 6.264 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.336 0.024 6.360 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.432 0.024 6.456 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.528 0.024 6.552 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.624 0.024 6.648 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.720 0.024 6.744 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.816 0.024 6.840 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.912 0.024 6.936 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.008 0.024 7.032 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.104 0.024 7.128 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.200 0.024 7.224 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.296 0.024 7.320 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.392 0.024 7.416 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.584 0.024 7.608 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.680 0.024 7.704 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.776 0.024 7.800 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.872 0.024 7.896 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.968 0.024 7.992 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.064 0.024 8.088 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.160 0.024 8.184 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.256 0.024 8.280 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.352 0.024 8.376 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.448 0.024 8.472 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.544 0.024 8.568 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.640 0.024 8.664 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.736 0.024 8.760 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.832 0.024 8.856 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.928 0.024 8.952 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.024 0.024 9.048 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.120 0.024 9.144 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.216 0.024 9.240 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.312 0.024 9.336 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.408 0.024 9.432 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.504 0.024 9.528 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.696 0.024 9.720 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.792 0.024 9.816 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.888 0.024 9.912 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.984 0.024 10.008 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.080 0.024 10.104 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.176 0.024 10.200 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.272 0.024 10.296 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.368 0.024 10.392 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.464 0.024 10.488 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.560 0.024 10.584 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.656 0.024 10.680 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.752 0.024 10.776 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.848 0.024 10.872 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.944 0.024 10.968 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.040 0.024 11.064 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.136 0.024 11.160 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.232 0.024 11.256 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END rd_out[117]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.840 0.024 15.864 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.936 0.024 15.960 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.032 0.024 16.056 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.128 0.024 16.152 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.224 0.024 16.248 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.320 0.024 16.344 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.416 0.024 16.440 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.512 0.024 16.536 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.608 0.024 16.632 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.704 0.024 16.728 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.800 0.024 16.824 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.896 0.024 16.920 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.992 0.024 17.016 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.088 0.024 17.112 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.184 0.024 17.208 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.280 0.024 17.304 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.376 0.024 17.400 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.472 0.024 17.496 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.568 0.024 17.592 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.664 0.024 17.688 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.760 0.024 17.784 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.856 0.024 17.880 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.952 0.024 17.976 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.048 0.024 18.072 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.144 0.024 18.168 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.240 0.024 18.264 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.336 0.024 18.360 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.432 0.024 18.456 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.528 0.024 18.552 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.624 0.024 18.648 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.720 0.024 18.744 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.816 0.024 18.840 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.912 0.024 18.936 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.008 0.024 19.032 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.104 0.024 19.128 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.200 0.024 19.224 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.296 0.024 19.320 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.392 0.024 19.416 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.488 0.024 19.512 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.584 0.024 19.608 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.680 0.024 19.704 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.776 0.024 19.800 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.872 0.024 19.896 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.968 0.024 19.992 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.064 0.024 20.088 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.160 0.024 20.184 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.256 0.024 20.280 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.352 0.024 20.376 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.448 0.024 20.472 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.544 0.024 20.568 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.640 0.024 20.664 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.736 0.024 20.760 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.832 0.024 20.856 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.928 0.024 20.952 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.024 0.024 21.048 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.120 0.024 21.144 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.216 0.024 21.240 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.312 0.024 21.336 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.408 0.024 21.432 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.504 0.024 21.528 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.600 0.024 21.624 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.696 0.024 21.720 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.792 0.024 21.816 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.888 0.024 21.912 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.984 0.024 22.008 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.080 0.024 22.104 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.176 0.024 22.200 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.272 0.024 22.296 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.368 0.024 22.392 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.464 0.024 22.488 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.560 0.024 22.584 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.656 0.024 22.680 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.752 0.024 22.776 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.848 0.024 22.872 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.944 0.024 22.968 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.040 0.024 23.064 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.136 0.024 23.160 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.232 0.024 23.256 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.328 0.024 23.352 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.424 0.024 23.448 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.520 0.024 23.544 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.616 0.024 23.640 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.712 0.024 23.736 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.808 0.024 23.832 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.904 0.024 23.928 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.000 0.024 24.024 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.096 0.024 24.120 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.192 0.024 24.216 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.288 0.024 24.312 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.384 0.024 24.408 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.480 0.024 24.504 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.576 0.024 24.600 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.672 0.024 24.696 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.768 0.024 24.792 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.864 0.024 24.888 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.960 0.024 24.984 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.056 0.024 25.080 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.152 0.024 25.176 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.248 0.024 25.272 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.344 0.024 25.368 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.440 0.024 25.464 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.536 0.024 25.560 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.632 0.024 25.656 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.728 0.024 25.752 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.824 0.024 25.848 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.920 0.024 25.944 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.016 0.024 26.040 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.112 0.024 26.136 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.208 0.024 26.232 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.304 0.024 26.328 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.400 0.024 26.424 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.496 0.024 26.520 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.592 0.024 26.616 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.688 0.024 26.712 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.784 0.024 26.808 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.880 0.024 26.904 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.976 0.024 27.000 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.072 0.024 27.096 ;
    END
  END wd_in[117]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.584 0.024 31.608 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.680 0.024 31.704 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.776 0.024 31.800 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.872 0.024 31.896 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.968 0.024 31.992 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.064 0.024 32.088 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.160 0.024 32.184 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.256 0.024 32.280 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.768 0.024 36.792 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.864 0.024 36.888 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.960 0.024 36.984 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 15.294 0.144 ;
      RECT 0.096 1.584 15.294 1.680 ;
      RECT 0.096 3.120 15.294 3.216 ;
      RECT 0.096 4.656 15.294 4.752 ;
      RECT 0.096 6.192 15.294 6.288 ;
      RECT 0.096 7.728 15.294 7.824 ;
      RECT 0.096 9.264 15.294 9.360 ;
      RECT 0.096 10.800 15.294 10.896 ;
      RECT 0.096 12.336 15.294 12.432 ;
      RECT 0.096 13.872 15.294 13.968 ;
      RECT 0.096 15.408 15.294 15.504 ;
      RECT 0.096 16.944 15.294 17.040 ;
      RECT 0.096 18.480 15.294 18.576 ;
      RECT 0.096 20.016 15.294 20.112 ;
      RECT 0.096 21.552 15.294 21.648 ;
      RECT 0.096 23.088 15.294 23.184 ;
      RECT 0.096 24.624 15.294 24.720 ;
      RECT 0.096 26.160 15.294 26.256 ;
      RECT 0.096 27.696 15.294 27.792 ;
      RECT 0.096 29.232 15.294 29.328 ;
      RECT 0.096 30.768 15.294 30.864 ;
      RECT 0.096 32.304 15.294 32.400 ;
      RECT 0.096 33.840 15.294 33.936 ;
      RECT 0.096 35.376 15.294 35.472 ;
      RECT 0.096 36.912 15.294 37.008 ;
      RECT 0.096 38.448 15.294 38.544 ;
      RECT 0.096 39.984 15.294 40.080 ;
      RECT 0.096 41.520 15.294 41.616 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 15.294 0.912 ;
      RECT 0.096 2.352 15.294 2.448 ;
      RECT 0.096 3.888 15.294 3.984 ;
      RECT 0.096 5.424 15.294 5.520 ;
      RECT 0.096 6.960 15.294 7.056 ;
      RECT 0.096 8.496 15.294 8.592 ;
      RECT 0.096 10.032 15.294 10.128 ;
      RECT 0.096 11.568 15.294 11.664 ;
      RECT 0.096 13.104 15.294 13.200 ;
      RECT 0.096 14.640 15.294 14.736 ;
      RECT 0.096 16.176 15.294 16.272 ;
      RECT 0.096 17.712 15.294 17.808 ;
      RECT 0.096 19.248 15.294 19.344 ;
      RECT 0.096 20.784 15.294 20.880 ;
      RECT 0.096 22.320 15.294 22.416 ;
      RECT 0.096 23.856 15.294 23.952 ;
      RECT 0.096 25.392 15.294 25.488 ;
      RECT 0.096 26.928 15.294 27.024 ;
      RECT 0.096 28.464 15.294 28.560 ;
      RECT 0.096 30.000 15.294 30.096 ;
      RECT 0.096 31.536 15.294 31.632 ;
      RECT 0.096 33.072 15.294 33.168 ;
      RECT 0.096 34.608 15.294 34.704 ;
      RECT 0.096 36.144 15.294 36.240 ;
      RECT 0.096 37.680 15.294 37.776 ;
      RECT 0.096 39.216 15.294 39.312 ;
      RECT 0.096 40.752 15.294 40.848 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 15.390 42.000 ;
    LAYER M2 ;
    RECT 0 0 15.390 42.000 ;
    LAYER M3 ;
    RECT 0 0 15.390 42.000 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 42.000 ;
    RECT 15.294 0 15.390 42.000 ;
    RECT 0.096 0.000 15.294 0.048 ;
    RECT 0.096 0.144 15.294 0.816 ;
    RECT 0.096 0.912 15.294 1.584 ;
    RECT 0.096 1.680 15.294 2.352 ;
    RECT 0.096 2.448 15.294 3.120 ;
    RECT 0.096 3.216 15.294 3.888 ;
    RECT 0.096 3.984 15.294 4.656 ;
    RECT 0.096 4.752 15.294 5.424 ;
    RECT 0.096 5.520 15.294 6.192 ;
    RECT 0.096 6.288 15.294 6.960 ;
    RECT 0.096 7.056 15.294 7.728 ;
    RECT 0.096 7.824 15.294 8.496 ;
    RECT 0.096 8.592 15.294 9.264 ;
    RECT 0.096 9.360 15.294 10.032 ;
    RECT 0.096 10.128 15.294 10.800 ;
    RECT 0.096 10.896 15.294 11.568 ;
    RECT 0.096 11.664 15.294 12.336 ;
    RECT 0.096 12.432 15.294 13.104 ;
    RECT 0.096 13.200 15.294 13.872 ;
    RECT 0.096 13.968 15.294 14.640 ;
    RECT 0.096 14.736 15.294 15.408 ;
    RECT 0.096 15.504 15.294 16.176 ;
    RECT 0.096 16.272 15.294 16.944 ;
    RECT 0.096 17.040 15.294 17.712 ;
    RECT 0.096 17.808 15.294 18.480 ;
    RECT 0.096 18.576 15.294 19.248 ;
    RECT 0.096 19.344 15.294 20.016 ;
    RECT 0.096 20.112 15.294 20.784 ;
    RECT 0.096 20.880 15.294 21.552 ;
    RECT 0.096 21.648 15.294 22.320 ;
    RECT 0.096 22.416 15.294 23.088 ;
    RECT 0.096 23.184 15.294 23.856 ;
    RECT 0.096 23.952 15.294 24.624 ;
    RECT 0.096 24.720 15.294 25.392 ;
    RECT 0.096 25.488 15.294 26.160 ;
    RECT 0.096 26.256 15.294 26.928 ;
    RECT 0.096 27.024 15.294 27.696 ;
    RECT 0.096 27.792 15.294 28.464 ;
    RECT 0.096 28.560 15.294 29.232 ;
    RECT 0.096 29.328 15.294 30.000 ;
    RECT 0.096 30.096 15.294 30.768 ;
    RECT 0.096 30.864 15.294 31.536 ;
    RECT 0.096 31.632 15.294 32.304 ;
    RECT 0.096 32.400 15.294 33.072 ;
    RECT 0.096 33.168 15.294 33.840 ;
    RECT 0.096 33.936 15.294 34.608 ;
    RECT 0.096 34.704 15.294 35.376 ;
    RECT 0.096 35.472 15.294 36.144 ;
    RECT 0.096 36.240 15.294 36.912 ;
    RECT 0.096 37.008 15.294 37.680 ;
    RECT 0.096 37.776 15.294 38.448 ;
    RECT 0.096 38.544 15.294 39.216 ;
    RECT 0.096 39.312 15.294 39.984 ;
    RECT 0.096 40.080 15.294 40.752 ;
    RECT 0.096 40.848 15.294 41.520 ;
    RECT 0.096 41.616 15.294 42.000 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 0.192 ;
    RECT 0 0.216 0.024 0.288 ;
    RECT 0 0.312 0.024 0.384 ;
    RECT 0 0.408 0.024 0.480 ;
    RECT 0 0.504 0.024 0.576 ;
    RECT 0 0.600 0.024 0.672 ;
    RECT 0 0.696 0.024 0.768 ;
    RECT 0 0.792 0.024 0.864 ;
    RECT 0 0.888 0.024 0.960 ;
    RECT 0 0.984 0.024 1.056 ;
    RECT 0 1.080 0.024 1.152 ;
    RECT 0 1.176 0.024 1.248 ;
    RECT 0 1.272 0.024 1.344 ;
    RECT 0 1.368 0.024 1.440 ;
    RECT 0 1.464 0.024 1.536 ;
    RECT 0 1.560 0.024 1.632 ;
    RECT 0 1.656 0.024 1.728 ;
    RECT 0 1.752 0.024 1.824 ;
    RECT 0 1.848 0.024 1.920 ;
    RECT 0 1.944 0.024 2.016 ;
    RECT 0 2.040 0.024 2.112 ;
    RECT 0 2.136 0.024 2.208 ;
    RECT 0 2.232 0.024 2.304 ;
    RECT 0 2.328 0.024 2.400 ;
    RECT 0 2.424 0.024 2.496 ;
    RECT 0 2.520 0.024 2.592 ;
    RECT 0 2.616 0.024 2.688 ;
    RECT 0 2.712 0.024 2.784 ;
    RECT 0 2.808 0.024 2.880 ;
    RECT 0 2.904 0.024 2.976 ;
    RECT 0 3.000 0.024 3.072 ;
    RECT 0 3.096 0.024 3.168 ;
    RECT 0 3.192 0.024 3.264 ;
    RECT 0 3.288 0.024 3.360 ;
    RECT 0 3.384 0.024 3.456 ;
    RECT 0 3.480 0.024 3.552 ;
    RECT 0 3.576 0.024 3.648 ;
    RECT 0 3.672 0.024 3.744 ;
    RECT 0 3.768 0.024 3.840 ;
    RECT 0 3.864 0.024 3.936 ;
    RECT 0 3.960 0.024 4.032 ;
    RECT 0 4.056 0.024 4.128 ;
    RECT 0 4.152 0.024 4.224 ;
    RECT 0 4.248 0.024 4.320 ;
    RECT 0 4.344 0.024 4.416 ;
    RECT 0 4.440 0.024 4.512 ;
    RECT 0 4.536 0.024 4.608 ;
    RECT 0 4.632 0.024 4.704 ;
    RECT 0 4.728 0.024 4.800 ;
    RECT 0 4.824 0.024 4.896 ;
    RECT 0 4.920 0.024 4.992 ;
    RECT 0 5.016 0.024 5.088 ;
    RECT 0 5.112 0.024 5.184 ;
    RECT 0 5.208 0.024 5.280 ;
    RECT 0 5.304 0.024 5.376 ;
    RECT 0 5.400 0.024 5.472 ;
    RECT 0 5.496 0.024 5.568 ;
    RECT 0 5.592 0.024 5.664 ;
    RECT 0 5.688 0.024 5.760 ;
    RECT 0 5.784 0.024 5.856 ;
    RECT 0 5.880 0.024 5.952 ;
    RECT 0 5.976 0.024 6.048 ;
    RECT 0 6.072 0.024 6.144 ;
    RECT 0 6.168 0.024 6.240 ;
    RECT 0 6.264 0.024 6.336 ;
    RECT 0 6.360 0.024 6.432 ;
    RECT 0 6.456 0.024 6.528 ;
    RECT 0 6.552 0.024 6.624 ;
    RECT 0 6.648 0.024 6.720 ;
    RECT 0 6.744 0.024 6.816 ;
    RECT 0 6.840 0.024 6.912 ;
    RECT 0 6.936 0.024 7.008 ;
    RECT 0 7.032 0.024 7.104 ;
    RECT 0 7.128 0.024 7.200 ;
    RECT 0 7.224 0.024 7.296 ;
    RECT 0 7.320 0.024 7.392 ;
    RECT 0 7.416 0.024 7.488 ;
    RECT 0 7.512 0.024 7.584 ;
    RECT 0 7.608 0.024 7.680 ;
    RECT 0 7.704 0.024 7.776 ;
    RECT 0 7.800 0.024 7.872 ;
    RECT 0 7.896 0.024 7.968 ;
    RECT 0 7.992 0.024 8.064 ;
    RECT 0 8.088 0.024 8.160 ;
    RECT 0 8.184 0.024 8.256 ;
    RECT 0 8.280 0.024 8.352 ;
    RECT 0 8.376 0.024 8.448 ;
    RECT 0 8.472 0.024 8.544 ;
    RECT 0 8.568 0.024 8.640 ;
    RECT 0 8.664 0.024 8.736 ;
    RECT 0 8.760 0.024 8.832 ;
    RECT 0 8.856 0.024 8.928 ;
    RECT 0 8.952 0.024 9.024 ;
    RECT 0 9.048 0.024 9.120 ;
    RECT 0 9.144 0.024 9.216 ;
    RECT 0 9.240 0.024 9.312 ;
    RECT 0 9.336 0.024 9.408 ;
    RECT 0 9.432 0.024 9.504 ;
    RECT 0 9.528 0.024 9.600 ;
    RECT 0 9.624 0.024 9.696 ;
    RECT 0 9.720 0.024 9.792 ;
    RECT 0 9.816 0.024 9.888 ;
    RECT 0 9.912 0.024 9.984 ;
    RECT 0 10.008 0.024 10.080 ;
    RECT 0 10.104 0.024 10.176 ;
    RECT 0 10.200 0.024 10.272 ;
    RECT 0 10.296 0.024 10.368 ;
    RECT 0 10.392 0.024 10.464 ;
    RECT 0 10.488 0.024 10.560 ;
    RECT 0 10.584 0.024 10.656 ;
    RECT 0 10.680 0.024 10.752 ;
    RECT 0 10.776 0.024 10.848 ;
    RECT 0 10.872 0.024 10.944 ;
    RECT 0 10.968 0.024 11.040 ;
    RECT 0 11.064 0.024 11.136 ;
    RECT 0 11.160 0.024 11.232 ;
    RECT 0 11.256 0.024 11.328 ;
    RECT 0 11.352 0.024 15.840 ;
    RECT 0 15.864 0.024 15.936 ;
    RECT 0 15.960 0.024 16.032 ;
    RECT 0 16.056 0.024 16.128 ;
    RECT 0 16.152 0.024 16.224 ;
    RECT 0 16.248 0.024 16.320 ;
    RECT 0 16.344 0.024 16.416 ;
    RECT 0 16.440 0.024 16.512 ;
    RECT 0 16.536 0.024 16.608 ;
    RECT 0 16.632 0.024 16.704 ;
    RECT 0 16.728 0.024 16.800 ;
    RECT 0 16.824 0.024 16.896 ;
    RECT 0 16.920 0.024 16.992 ;
    RECT 0 17.016 0.024 17.088 ;
    RECT 0 17.112 0.024 17.184 ;
    RECT 0 17.208 0.024 17.280 ;
    RECT 0 17.304 0.024 17.376 ;
    RECT 0 17.400 0.024 17.472 ;
    RECT 0 17.496 0.024 17.568 ;
    RECT 0 17.592 0.024 17.664 ;
    RECT 0 17.688 0.024 17.760 ;
    RECT 0 17.784 0.024 17.856 ;
    RECT 0 17.880 0.024 17.952 ;
    RECT 0 17.976 0.024 18.048 ;
    RECT 0 18.072 0.024 18.144 ;
    RECT 0 18.168 0.024 18.240 ;
    RECT 0 18.264 0.024 18.336 ;
    RECT 0 18.360 0.024 18.432 ;
    RECT 0 18.456 0.024 18.528 ;
    RECT 0 18.552 0.024 18.624 ;
    RECT 0 18.648 0.024 18.720 ;
    RECT 0 18.744 0.024 18.816 ;
    RECT 0 18.840 0.024 18.912 ;
    RECT 0 18.936 0.024 19.008 ;
    RECT 0 19.032 0.024 19.104 ;
    RECT 0 19.128 0.024 19.200 ;
    RECT 0 19.224 0.024 19.296 ;
    RECT 0 19.320 0.024 19.392 ;
    RECT 0 19.416 0.024 19.488 ;
    RECT 0 19.512 0.024 19.584 ;
    RECT 0 19.608 0.024 19.680 ;
    RECT 0 19.704 0.024 19.776 ;
    RECT 0 19.800 0.024 19.872 ;
    RECT 0 19.896 0.024 19.968 ;
    RECT 0 19.992 0.024 20.064 ;
    RECT 0 20.088 0.024 20.160 ;
    RECT 0 20.184 0.024 20.256 ;
    RECT 0 20.280 0.024 20.352 ;
    RECT 0 20.376 0.024 20.448 ;
    RECT 0 20.472 0.024 20.544 ;
    RECT 0 20.568 0.024 20.640 ;
    RECT 0 20.664 0.024 20.736 ;
    RECT 0 20.760 0.024 20.832 ;
    RECT 0 20.856 0.024 20.928 ;
    RECT 0 20.952 0.024 21.024 ;
    RECT 0 21.048 0.024 21.120 ;
    RECT 0 21.144 0.024 21.216 ;
    RECT 0 21.240 0.024 21.312 ;
    RECT 0 21.336 0.024 21.408 ;
    RECT 0 21.432 0.024 21.504 ;
    RECT 0 21.528 0.024 21.600 ;
    RECT 0 21.624 0.024 21.696 ;
    RECT 0 21.720 0.024 21.792 ;
    RECT 0 21.816 0.024 21.888 ;
    RECT 0 21.912 0.024 21.984 ;
    RECT 0 22.008 0.024 22.080 ;
    RECT 0 22.104 0.024 22.176 ;
    RECT 0 22.200 0.024 22.272 ;
    RECT 0 22.296 0.024 22.368 ;
    RECT 0 22.392 0.024 22.464 ;
    RECT 0 22.488 0.024 22.560 ;
    RECT 0 22.584 0.024 22.656 ;
    RECT 0 22.680 0.024 22.752 ;
    RECT 0 22.776 0.024 22.848 ;
    RECT 0 22.872 0.024 22.944 ;
    RECT 0 22.968 0.024 23.040 ;
    RECT 0 23.064 0.024 23.136 ;
    RECT 0 23.160 0.024 23.232 ;
    RECT 0 23.256 0.024 23.328 ;
    RECT 0 23.352 0.024 23.424 ;
    RECT 0 23.448 0.024 23.520 ;
    RECT 0 23.544 0.024 23.616 ;
    RECT 0 23.640 0.024 23.712 ;
    RECT 0 23.736 0.024 23.808 ;
    RECT 0 23.832 0.024 23.904 ;
    RECT 0 23.928 0.024 24.000 ;
    RECT 0 24.024 0.024 24.096 ;
    RECT 0 24.120 0.024 24.192 ;
    RECT 0 24.216 0.024 24.288 ;
    RECT 0 24.312 0.024 24.384 ;
    RECT 0 24.408 0.024 24.480 ;
    RECT 0 24.504 0.024 24.576 ;
    RECT 0 24.600 0.024 24.672 ;
    RECT 0 24.696 0.024 24.768 ;
    RECT 0 24.792 0.024 24.864 ;
    RECT 0 24.888 0.024 24.960 ;
    RECT 0 24.984 0.024 25.056 ;
    RECT 0 25.080 0.024 25.152 ;
    RECT 0 25.176 0.024 25.248 ;
    RECT 0 25.272 0.024 25.344 ;
    RECT 0 25.368 0.024 25.440 ;
    RECT 0 25.464 0.024 25.536 ;
    RECT 0 25.560 0.024 25.632 ;
    RECT 0 25.656 0.024 25.728 ;
    RECT 0 25.752 0.024 25.824 ;
    RECT 0 25.848 0.024 25.920 ;
    RECT 0 25.944 0.024 26.016 ;
    RECT 0 26.040 0.024 26.112 ;
    RECT 0 26.136 0.024 26.208 ;
    RECT 0 26.232 0.024 26.304 ;
    RECT 0 26.328 0.024 26.400 ;
    RECT 0 26.424 0.024 26.496 ;
    RECT 0 26.520 0.024 26.592 ;
    RECT 0 26.616 0.024 26.688 ;
    RECT 0 26.712 0.024 26.784 ;
    RECT 0 26.808 0.024 26.880 ;
    RECT 0 26.904 0.024 26.976 ;
    RECT 0 27.000 0.024 27.072 ;
    RECT 0 27.096 0.024 31.584 ;
    RECT 0 31.608 0.024 31.680 ;
    RECT 0 31.704 0.024 31.776 ;
    RECT 0 31.800 0.024 31.872 ;
    RECT 0 31.896 0.024 31.968 ;
    RECT 0 31.992 0.024 32.064 ;
    RECT 0 32.088 0.024 32.160 ;
    RECT 0 32.184 0.024 32.256 ;
    RECT 0 32.280 0.024 32.352 ;
    RECT 0 32.376 0.024 32.448 ;
    RECT 0 32.472 0.024 32.544 ;
    RECT 0 32.568 0.024 32.640 ;
    RECT 0 32.664 0.024 32.736 ;
    RECT 0 32.760 0.024 32.832 ;
    RECT 0 32.856 0.024 32.928 ;
    RECT 0 32.952 0.024 33.024 ;
    RECT 0 33.048 0.024 33.120 ;
    RECT 0 33.144 0.024 33.216 ;
    RECT 0 33.240 0.024 33.312 ;
    RECT 0 33.336 0.024 33.408 ;
    RECT 0 33.432 0.024 33.504 ;
    RECT 0 33.528 0.024 33.600 ;
    RECT 0 33.624 0.024 33.696 ;
    RECT 0 33.720 0.024 33.792 ;
    RECT 0 33.816 0.024 33.888 ;
    RECT 0 33.912 0.024 33.984 ;
    RECT 0 34.008 0.024 34.080 ;
    RECT 0 34.104 0.024 34.176 ;
    RECT 0 34.200 0.024 34.272 ;
    RECT 0 34.296 0.024 34.368 ;
    RECT 0 34.392 0.024 34.464 ;
    RECT 0 34.488 0.024 34.560 ;
    RECT 0 34.584 0.024 34.656 ;
    RECT 0 34.680 0.024 34.752 ;
    RECT 0 34.776 0.024 34.848 ;
    RECT 0 34.872 0.024 34.944 ;
    RECT 0 34.968 0.024 35.040 ;
    RECT 0 35.064 0.024 35.136 ;
    RECT 0 35.160 0.024 35.232 ;
    RECT 0 35.256 0.024 35.328 ;
    RECT 0 35.352 0.024 35.424 ;
    RECT 0 35.448 0.024 35.520 ;
    RECT 0 35.544 0.024 35.616 ;
    RECT 0 35.640 0.024 35.712 ;
    RECT 0 35.736 0.024 35.808 ;
    RECT 0 35.832 0.024 35.904 ;
    RECT 0 35.928 0.024 36.000 ;
    RECT 0 36.024 0.024 36.096 ;
    RECT 0 36.120 0.024 36.192 ;
    RECT 0 36.216 0.024 36.288 ;
    RECT 0 36.312 0.024 36.384 ;
    RECT 0 36.408 0.024 36.480 ;
    RECT 0 36.504 0.024 36.576 ;
    RECT 0 36.600 0.024 36.672 ;
    RECT 0 36.696 0.024 36.768 ;
    RECT 0 36.792 0.024 36.864 ;
    RECT 0 36.888 0.024 36.960 ;
    RECT 0 36.984 0.024 37.056 ;
    RECT 0 37.080 0.024 37.152 ;
    RECT 0 37.176 0.024 37.248 ;
    RECT 0 37.272 0.024 37.344 ;
    RECT 0 37.368 0.024 37.440 ;
    RECT 0 37.464 0.024 37.536 ;
    RECT 0 37.560 0.024 37.632 ;
    RECT 0 37.656 0.024 37.728 ;
    RECT 0 37.752 0.024 37.824 ;
    RECT 0 37.848 0.024 37.920 ;
    RECT 0 37.944 0.024 38.016 ;
    RECT 0 38.040 0.024 38.112 ;
    RECT 0 38.136 0.024 38.208 ;
    RECT 0 38.232 0.024 38.304 ;
    RECT 0 38.328 0.024 38.400 ;
    RECT 0 38.424 0.024 38.496 ;
    RECT 0 38.520 0.024 38.592 ;
    RECT 0 38.616 0.024 38.688 ;
    RECT 0 38.712 0.024 38.784 ;
    RECT 0 38.808 0.024 38.880 ;
    RECT 0 38.904 0.024 38.976 ;
    RECT 0 39.000 0.024 39.072 ;
    RECT 0 39.096 0.024 39.168 ;
    RECT 0 39.192 0.024 39.264 ;
    RECT 0 39.288 0.024 39.360 ;
    RECT 0 39.384 0.024 39.456 ;
    RECT 0 39.480 0.024 39.552 ;
    RECT 0 39.576 0.024 39.648 ;
    RECT 0 39.672 0.024 39.744 ;
    RECT 0 39.768 0.024 39.840 ;
    RECT 0 39.864 0.024 39.936 ;
    RECT 0 39.960 0.024 40.032 ;
    RECT 0 40.056 0.024 40.128 ;
    RECT 0 40.152 0.024 40.224 ;
    RECT 0 40.248 0.024 40.320 ;
    RECT 0 40.344 0.024 40.416 ;
    RECT 0 40.440 0.024 40.512 ;
    RECT 0 40.536 0.024 40.608 ;
    RECT 0 40.632 0.024 40.704 ;
    RECT 0 40.728 0.024 40.800 ;
    RECT 0 40.824 0.024 40.896 ;
    RECT 0 40.920 0.024 40.992 ;
    RECT 0 41.016 0.024 41.088 ;
    RECT 0 41.112 0.024 41.184 ;
    RECT 0 41.208 0.024 41.280 ;
    RECT 0 41.304 0.024 41.376 ;
    RECT 0 41.400 0.024 41.472 ;
    RECT 0 41.496 0.024 41.568 ;
    RECT 0 41.592 0.024 41.664 ;
    RECT 0 41.688 0.024 41.760 ;
    RECT 0 41.784 0.024 41.856 ;
    RECT 0 41.880 0.024 41.952 ;
    RECT 0 41.976 0.024 42.048 ;
    RECT 0 42.072 0.024 42.144 ;
    RECT 0 42.168 0.024 42.240 ;
    RECT 0 42.264 0.024 42.336 ;
    RECT 0 42.360 0.024 42.432 ;
    RECT 0 42.456 0.024 42.528 ;
    RECT 0 42.552 0.024 42.624 ;
    RECT 0 42.648 0.024 42.720 ;
    RECT 0 42.744 0.024 42.816 ;
    RECT 0 42.840 0.024 47.328 ;
    RECT 0 47.352 0.024 47.424 ;
    RECT 0 47.448 0.024 47.520 ;
    RECT 0 47.544 0.024 47.616 ;
    RECT 0 47.640 0.024 47.712 ;
    RECT 0 47.736 0.024 47.808 ;
    RECT 0 47.832 0.024 47.904 ;
    RECT 0 47.928 0.024 48.000 ;
    RECT 0 48.024 0.024 52.512 ;
    RECT 0 52.536 0.024 52.608 ;
    RECT 0 52.632 0.024 52.704 ;
    RECT 0 52.728 0.024 42.000 ;
    LAYER OVERLAP ;
    RECT 0 0 15.390 42.000 ;
  END
END fakeram7_160x118

END LIBRARY
