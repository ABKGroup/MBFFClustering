VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE asap7sc7p5t_R8
  CLASS CORE ;
  SIZE 0.054 BY 2.16 ;
  SYMMETRY Y ;
END asap7sc7p5t_R8

MACRO DFFHQNV8H2Xx2_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0.0 0.0 ;
  FOREIGN DFFHQNV8H2Xx2_ASAP7_75t_SL 0.0 0.0 ;
  SIZE 2.268 BY 2.16 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_R8 ;
    PIN VDD
      USE POWER ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 0.261 1.134 0.279 ;
          RECT 1.134 0.261 2.268 0.279 ;
          RECT 0.0 0.801 1.134 0.819 ;
          RECT 1.134 0.801 2.268 0.819 ;
          RECT 0.0 1.341 1.134 1.359 ;
          RECT 1.134 1.341 2.268 1.359 ;
          RECT 0.0 1.881 1.134 1.899 ;
          RECT 1.134 1.881 2.268 1.899 ;
      END
    END VDD
    PIN VSS
      USE GROUND ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 -0.009 1.134 0.009 ;
          RECT 1.134 -0.009 2.268 0.009 ;
          RECT 0.0 0.549 1.134 0.531 ;
          RECT 1.134 0.549 2.268 0.531 ;
          RECT 0.0 1.089 1.134 1.071 ;
          RECT 1.134 1.089 2.268 1.071 ;
          RECT 0.0 1.629 1.134 1.611 ;
          RECT 1.134 1.629 2.268 1.611 ;
          RECT 0.0 2.169 1.134 2.151 ;
          RECT 1.134 2.169 2.268 2.151 ;
      END
    END VSS
    PIN CLK
      USE CLOCK ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.099 0.164 0.117 0.236 ;
          RECT 0.072 0.07 0.117 0.106 ;
          RECT 0.099 0.034 0.117 0.106 ;
          RECT 0.072 0.164 0.117 0.2 ;
          RECT 0.072 0.07 0.09 0.2 ;
          RECT 1.233 0.164 1.251 0.236 ;
          RECT 1.206 0.07 1.251 0.106 ;
          RECT 1.233 0.034 1.251 0.106 ;
          RECT 1.206 0.164 1.251 0.2 ;
          RECT 1.206 0.07 1.224 0.2 ;
          RECT 0.099 0.376 0.117 0.304 ;
          RECT 0.072 0.47 0.117 0.434 ;
          RECT 0.099 0.506 0.117 0.434 ;
          RECT 0.072 0.376 0.117 0.34 ;
          RECT 0.072 0.47 0.09 0.34 ;
          RECT 1.233 0.376 1.251 0.304 ;
          RECT 1.206 0.47 1.251 0.434 ;
          RECT 1.233 0.506 1.251 0.434 ;
          RECT 1.206 0.376 1.251 0.34 ;
          RECT 1.206 0.47 1.224 0.34 ;
          RECT 0.099 0.704 0.117 0.776 ;
          RECT 0.072 0.61 0.117 0.646 ;
          RECT 0.099 0.574 0.117 0.646 ;
          RECT 0.072 0.704 0.117 0.74 ;
          RECT 0.072 0.61 0.09 0.74 ;
          RECT 1.233 0.704 1.251 0.776 ;
          RECT 1.206 0.61 1.251 0.646 ;
          RECT 1.233 0.574 1.251 0.646 ;
          RECT 1.206 0.704 1.251 0.74 ;
          RECT 1.206 0.61 1.224 0.74 ;
          RECT 0.099 0.916 0.117 0.844 ;
          RECT 0.072 1.01 0.117 0.974 ;
          RECT 0.099 1.046 0.117 0.974 ;
          RECT 0.072 0.916 0.117 0.88 ;
          RECT 0.072 1.01 0.09 0.88 ;
          RECT 1.233 0.916 1.251 0.844 ;
          RECT 1.206 1.01 1.251 0.974 ;
          RECT 1.233 1.046 1.251 0.974 ;
          RECT 1.206 0.916 1.251 0.88 ;
          RECT 1.206 1.01 1.224 0.88 ;
          RECT 0.099 1.244 0.117 1.316 ;
          RECT 0.072 1.15 0.117 1.186 ;
          RECT 0.099 1.114 0.117 1.186 ;
          RECT 0.072 1.244 0.117 1.28 ;
          RECT 0.072 1.15 0.09 1.28 ;
          RECT 1.233 1.244 1.251 1.316 ;
          RECT 1.206 1.15 1.251 1.186 ;
          RECT 1.233 1.114 1.251 1.186 ;
          RECT 1.206 1.244 1.251 1.28 ;
          RECT 1.206 1.15 1.224 1.28 ;
          RECT 0.099 1.456 0.117 1.384 ;
          RECT 0.072 1.55 0.117 1.514 ;
          RECT 0.099 1.586 0.117 1.514 ;
          RECT 0.072 1.456 0.117 1.42 ;
          RECT 0.072 1.55 0.09 1.42 ;
          RECT 1.233 1.456 1.251 1.384 ;
          RECT 1.206 1.55 1.251 1.514 ;
          RECT 1.233 1.586 1.251 1.514 ;
          RECT 1.206 1.456 1.251 1.42 ;
          RECT 1.206 1.55 1.224 1.42 ;
          RECT 0.099 1.784 0.117 1.856 ;
          RECT 0.072 1.69 0.117 1.726 ;
          RECT 0.099 1.654 0.117 1.726 ;
          RECT 0.072 1.784 0.117 1.82 ;
          RECT 0.072 1.69 0.09 1.82 ;
          RECT 1.233 1.784 1.251 1.856 ;
          RECT 1.206 1.69 1.251 1.726 ;
          RECT 1.233 1.654 1.251 1.726 ;
          RECT 1.206 1.784 1.251 1.82 ;
          RECT 1.206 1.69 1.224 1.82 ;
          RECT 0.099 1.996 0.117 1.924 ;
          RECT 0.072 2.09 0.117 2.054 ;
          RECT 0.099 2.126 0.117 2.054 ;
          RECT 0.072 1.996 0.117 1.96 ;
          RECT 0.072 2.09 0.09 1.96 ;
          RECT 1.233 1.996 1.251 1.924 ;
          RECT 1.206 2.09 1.251 2.054 ;
          RECT 1.233 2.126 1.251 2.054 ;
          RECT 1.206 1.996 1.251 1.96 ;
          RECT 1.206 2.09 1.224 1.96 ;
        LAYER M2 ;
          RECT 0.072 0.072 1.35 0.09 ;
          RECT 0.072 0.45 1.35 0.468 ;
          RECT 0.072 0.612 1.35 0.63 ;
          RECT 0.072 0.99 1.35 1.008 ;
          RECT 0.072 1.152 1.35 1.17 ;
          RECT 0.072 1.53 1.35 1.548 ;
          RECT 0.072 1.692 1.35 1.71 ;
          RECT 0.072 2.07 1.35 2.088 ;
        LAYER V1 ;
          RECT 0.099 0.072 0.117 0.09 ;
          RECT 1.233 0.072 1.251 0.09 ;
          RECT 0.099 0.45 0.117 0.468 ;
          RECT 1.233 0.45 1.251 0.468 ;
          RECT 0.099 0.612 0.117 0.63 ;
          RECT 1.233 0.612 1.251 0.63 ;
          RECT 0.099 0.99 0.117 1.008 ;
          RECT 1.233 0.99 1.251 1.008 ;
          RECT 0.099 1.152 0.117 1.17 ;
          RECT 1.233 1.152 1.251 1.17 ;
          RECT 0.099 1.53 0.117 1.548 ;
          RECT 1.233 1.53 1.251 1.548 ;
          RECT 0.099 1.692 0.117 1.71 ;
          RECT 1.233 1.692 1.251 1.71 ;
          RECT 0.099 2.07 0.117 2.088 ;
          RECT 1.233 2.07 1.251 2.088 ;
        LAYER M3 ;
          RECT 0.171 0.054 0.189 2.106 ;
        LAYER V2 ;
          RECT 0.171 0.072 0.189 0.09 ;
          RECT 0.171 0.45 0.189 0.468 ;
          RECT 0.171 0.612 0.189 0.63 ;
          RECT 0.171 0.99 0.189 1.008 ;
          RECT 0.171 1.152 0.189 1.17 ;
          RECT 0.171 1.53 0.189 1.548 ;
          RECT 0.171 1.692 0.189 1.71 ;
          RECT 0.171 2.07 0.189 2.088 ;
      END
    END CLK
    PIN D0
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.126 0.29 0.144 ;
          RECT 0.234 0.225 0.271 0.243 ;
          RECT 0.234 0.027 0.271 0.045 ;
          RECT 0.234 0.027 0.252 0.243 ;
      END
    END D0
    PIN QN0
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.216 1.117 0.234 ;
          RECT 1.099 0.036 1.117 0.234 ;
          RECT 1.012 0.036 1.117 0.054 ;
      END
    END QN0
    PIN D1
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 0.126 1.424 0.144 ;
          RECT 1.368 0.225 1.405 0.243 ;
          RECT 1.368 0.027 1.405 0.045 ;
          RECT 1.368 0.027 1.386 0.243 ;
      END
    END D1
    PIN QN1
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 0.216 2.251 0.234 ;
          RECT 2.233 0.036 2.251 0.234 ;
          RECT 2.146 0.036 2.251 0.054 ;
      END
    END QN1
    PIN D2
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.414 0.29 0.396 ;
          RECT 0.234 0.315 0.271 0.297 ;
          RECT 0.234 0.513 0.271 0.495 ;
          RECT 0.234 0.513 0.252 0.297 ;
      END
    END D2
    PIN QN2
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.324 1.117 0.306 ;
          RECT 1.099 0.504 1.117 0.306 ;
          RECT 1.012 0.504 1.117 0.486 ;
      END
    END QN2
    PIN D3
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 0.414 1.424 0.396 ;
          RECT 1.368 0.315 1.405 0.297 ;
          RECT 1.368 0.513 1.405 0.495 ;
          RECT 1.368 0.513 1.386 0.297 ;
      END
    END D3
    PIN QN3
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 0.324 2.251 0.306 ;
          RECT 2.233 0.504 2.251 0.306 ;
          RECT 2.146 0.504 2.251 0.486 ;
      END
    END QN3
    PIN D4
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.666 0.29 0.684 ;
          RECT 0.234 0.765 0.271 0.783 ;
          RECT 0.234 0.567 0.271 0.585 ;
          RECT 0.234 0.567 0.252 0.783 ;
      END
    END D4
    PIN QN4
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.756 1.117 0.774 ;
          RECT 1.099 0.576 1.117 0.774 ;
          RECT 1.012 0.576 1.117 0.594 ;
      END
    END QN4
    PIN D5
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 0.666 1.424 0.684 ;
          RECT 1.368 0.765 1.405 0.783 ;
          RECT 1.368 0.567 1.405 0.585 ;
          RECT 1.368 0.567 1.386 0.783 ;
      END
    END D5
    PIN QN5
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 0.756 2.251 0.774 ;
          RECT 2.233 0.576 2.251 0.774 ;
          RECT 2.146 0.576 2.251 0.594 ;
      END
    END QN5
    PIN D6
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.954 0.29 0.936 ;
          RECT 0.234 0.855 0.271 0.837 ;
          RECT 0.234 1.053 0.271 1.035 ;
          RECT 0.234 1.053 0.252 0.837 ;
      END
    END D6
    PIN QN6
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.864 1.117 0.846 ;
          RECT 1.099 1.044 1.117 0.846 ;
          RECT 1.012 1.044 1.117 1.026 ;
      END
    END QN6
    PIN D7
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 0.954 1.424 0.936 ;
          RECT 1.368 0.855 1.405 0.837 ;
          RECT 1.368 1.053 1.405 1.035 ;
          RECT 1.368 1.053 1.386 0.837 ;
      END
    END D7
    PIN QN7
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 0.864 2.251 0.846 ;
          RECT 2.233 1.044 2.251 0.846 ;
          RECT 2.146 1.044 2.251 1.026 ;
      END
    END QN7
    PIN D8
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.206 0.29 1.224 ;
          RECT 0.234 1.305 0.271 1.323 ;
          RECT 0.234 1.107 0.271 1.125 ;
          RECT 0.234 1.107 0.252 1.323 ;
      END
    END D8
    PIN QN8
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.296 1.117 1.314 ;
          RECT 1.099 1.116 1.117 1.314 ;
          RECT 1.012 1.116 1.117 1.134 ;
      END
    END QN8
    PIN D9
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 1.206 1.424 1.224 ;
          RECT 1.368 1.305 1.405 1.323 ;
          RECT 1.368 1.107 1.405 1.125 ;
          RECT 1.368 1.107 1.386 1.323 ;
      END
    END D9
    PIN QN9
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 1.296 2.251 1.314 ;
          RECT 2.233 1.116 2.251 1.314 ;
          RECT 2.146 1.116 2.251 1.134 ;
      END
    END QN9
    PIN D10
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.494 0.29 1.476 ;
          RECT 0.234 1.395 0.271 1.377 ;
          RECT 0.234 1.593 0.271 1.575 ;
          RECT 0.234 1.593 0.252 1.377 ;
      END
    END D10
    PIN QN10
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.404 1.117 1.386 ;
          RECT 1.099 1.584 1.117 1.386 ;
          RECT 1.012 1.584 1.117 1.566 ;
      END
    END QN10
    PIN D11
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 1.494 1.424 1.476 ;
          RECT 1.368 1.395 1.405 1.377 ;
          RECT 1.368 1.593 1.405 1.575 ;
          RECT 1.368 1.593 1.386 1.377 ;
      END
    END D11
    PIN QN11
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 1.404 2.251 1.386 ;
          RECT 2.233 1.584 2.251 1.386 ;
          RECT 2.146 1.584 2.251 1.566 ;
      END
    END QN11
    PIN D12
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.746 0.29 1.764 ;
          RECT 0.234 1.845 0.271 1.863 ;
          RECT 0.234 1.647 0.271 1.665 ;
          RECT 0.234 1.647 0.252 1.863 ;
      END
    END D12
    PIN QN12
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.836 1.117 1.854 ;
          RECT 1.099 1.656 1.117 1.854 ;
          RECT 1.012 1.656 1.117 1.674 ;
      END
    END QN12
    PIN D13
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 1.746 1.424 1.764 ;
          RECT 1.368 1.845 1.405 1.863 ;
          RECT 1.368 1.647 1.405 1.665 ;
          RECT 1.368 1.647 1.386 1.863 ;
      END
    END D13
    PIN QN13
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 1.836 2.251 1.854 ;
          RECT 2.233 1.656 2.251 1.854 ;
          RECT 2.146 1.656 2.251 1.674 ;
      END
    END QN13
    PIN D14
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 2.034 0.29 2.016 ;
          RECT 0.234 1.935 0.271 1.917 ;
          RECT 0.234 2.133 0.271 2.115 ;
          RECT 0.234 2.133 0.252 1.917 ;
      END
    END D14
    PIN QN14
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.944 1.117 1.926 ;
          RECT 1.099 2.124 1.117 1.926 ;
          RECT 1.012 2.124 1.117 2.106 ;
      END
    END QN14
    PIN D15
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.368 2.034 1.424 2.016 ;
          RECT 1.368 1.935 1.405 1.917 ;
          RECT 1.368 2.133 1.405 2.115 ;
          RECT 1.368 2.133 1.386 1.917 ;
      END
    END D15
    PIN QN15
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.146 1.944 2.251 1.926 ;
          RECT 2.233 2.124 2.251 1.926 ;
          RECT 2.146 2.124 2.251 2.106 ;
      END
    END QN15
    OBS
      LAYER M1 ;
        RECT 0.85 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.774 0.027 0.792 0.119 ;
        RECT 0.774 0.027 0.954 0.045 ;
        RECT 0.688 0.224 0.738 0.242 ;
        RECT 0.72 0.027 0.738 0.242 ;
        RECT 0.72 0.153 0.9 0.171 ;
        RECT 0.882 0.117 0.9 0.171 ;
        RECT 0.828 0.117 0.846 0.171 ;
        RECT 0.634 0.027 0.738 0.045 ;
        RECT 0.576 0.225 0.63 0.243 ;
        RECT 0.612 0.081 0.63 0.243 ;
        RECT 0.496 0.081 0.63 0.099 ;
        RECT 0.585 0.045 0.603 0.099 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.45 0.122 0.576 0.14 ;
        RECT 0.418 0.027 0.468 0.045 ;
        RECT 0.315 0.126 0.333 0.203 ;
        RECT 0.315 0.126 0.367 0.144 ;
        RECT 0.148 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.148 0.027 0.198 0.045 ;
        RECT 0.009 0.225 0.068 0.243 ;
        RECT 0.009 0.027 0.027 0.243 ;
        RECT 0.009 0.144 0.047 0.162 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.99 0.09 1.008 0.167 ;
        RECT 0.666 0.101 0.684 0.167 ;
        RECT 0.504 0.165 0.522 0.203 ;
        RECT 0.396 0.106 0.414 0.167 ;
        RECT 0.142 0.106 0.16 0.167 ;
        RECT 1.984 0.225 2.088 0.243 ;
        RECT 2.07 0.027 2.088 0.243 ;
        RECT 1.908 0.027 1.926 0.119 ;
        RECT 1.908 0.027 2.088 0.045 ;
        RECT 1.822 0.224 1.872 0.242 ;
        RECT 1.854 0.027 1.872 0.242 ;
        RECT 1.854 0.153 2.034 0.171 ;
        RECT 2.016 0.117 2.034 0.171 ;
        RECT 1.962 0.117 1.98 0.171 ;
        RECT 1.768 0.027 1.872 0.045 ;
        RECT 1.71 0.225 1.764 0.243 ;
        RECT 1.746 0.081 1.764 0.243 ;
        RECT 1.63 0.081 1.764 0.099 ;
        RECT 1.719 0.045 1.737 0.099 ;
        RECT 1.498 0.225 1.602 0.243 ;
        RECT 1.584 0.027 1.602 0.243 ;
        RECT 1.584 0.122 1.71 0.14 ;
        RECT 1.552 0.027 1.602 0.045 ;
        RECT 1.449 0.126 1.467 0.203 ;
        RECT 1.449 0.126 1.501 0.144 ;
        RECT 1.282 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.282 0.027 1.332 0.045 ;
        RECT 1.143 0.225 1.202 0.243 ;
        RECT 1.143 0.027 1.161 0.243 ;
        RECT 1.143 0.144 1.181 0.162 ;
        RECT 1.143 0.027 1.202 0.045 ;
        RECT 2.124 0.09 2.142 0.167 ;
        RECT 1.8 0.101 1.818 0.167 ;
        RECT 1.638 0.165 1.656 0.203 ;
        RECT 1.53 0.106 1.548 0.167 ;
        RECT 1.276 0.106 1.294 0.167 ;
        RECT 0.85 0.315 0.954 0.297 ;
        RECT 0.936 0.513 0.954 0.297 ;
        RECT 0.774 0.513 0.792 0.421 ;
        RECT 0.774 0.513 0.954 0.495 ;
        RECT 0.688 0.316 0.738 0.298 ;
        RECT 0.72 0.513 0.738 0.298 ;
        RECT 0.72 0.387 0.9 0.369 ;
        RECT 0.882 0.423 0.9 0.369 ;
        RECT 0.828 0.423 0.846 0.369 ;
        RECT 0.634 0.513 0.738 0.495 ;
        RECT 0.576 0.315 0.63 0.297 ;
        RECT 0.612 0.459 0.63 0.297 ;
        RECT 0.496 0.459 0.63 0.441 ;
        RECT 0.585 0.495 0.603 0.441 ;
        RECT 0.364 0.315 0.468 0.297 ;
        RECT 0.45 0.513 0.468 0.297 ;
        RECT 0.45 0.418 0.576 0.4 ;
        RECT 0.418 0.513 0.468 0.495 ;
        RECT 0.315 0.414 0.333 0.337 ;
        RECT 0.315 0.414 0.367 0.396 ;
        RECT 0.148 0.315 0.198 0.297 ;
        RECT 0.18 0.513 0.198 0.297 ;
        RECT 0.148 0.513 0.198 0.495 ;
        RECT 0.009 0.315 0.068 0.297 ;
        RECT 0.009 0.513 0.027 0.297 ;
        RECT 0.009 0.396 0.047 0.378 ;
        RECT 0.009 0.513 0.068 0.495 ;
        RECT 0.99 0.45 1.008 0.373 ;
        RECT 0.666 0.439 0.684 0.373 ;
        RECT 0.504 0.375 0.522 0.337 ;
        RECT 0.396 0.434 0.414 0.373 ;
        RECT 0.142 0.434 0.16 0.373 ;
        RECT 1.984 0.315 2.088 0.297 ;
        RECT 2.07 0.513 2.088 0.297 ;
        RECT 1.908 0.513 1.926 0.421 ;
        RECT 1.908 0.513 2.088 0.495 ;
        RECT 1.822 0.316 1.872 0.298 ;
        RECT 1.854 0.513 1.872 0.298 ;
        RECT 1.854 0.387 2.034 0.369 ;
        RECT 2.016 0.423 2.034 0.369 ;
        RECT 1.962 0.423 1.98 0.369 ;
        RECT 1.768 0.513 1.872 0.495 ;
        RECT 1.71 0.315 1.764 0.297 ;
        RECT 1.746 0.459 1.764 0.297 ;
        RECT 1.63 0.459 1.764 0.441 ;
        RECT 1.719 0.495 1.737 0.441 ;
        RECT 1.498 0.315 1.602 0.297 ;
        RECT 1.584 0.513 1.602 0.297 ;
        RECT 1.584 0.418 1.71 0.4 ;
        RECT 1.552 0.513 1.602 0.495 ;
        RECT 1.449 0.414 1.467 0.337 ;
        RECT 1.449 0.414 1.501 0.396 ;
        RECT 1.282 0.315 1.332 0.297 ;
        RECT 1.314 0.513 1.332 0.297 ;
        RECT 1.282 0.513 1.332 0.495 ;
        RECT 1.143 0.315 1.202 0.297 ;
        RECT 1.143 0.513 1.161 0.297 ;
        RECT 1.143 0.396 1.181 0.378 ;
        RECT 1.143 0.513 1.202 0.495 ;
        RECT 2.124 0.45 2.142 0.373 ;
        RECT 1.8 0.439 1.818 0.373 ;
        RECT 1.638 0.375 1.656 0.337 ;
        RECT 1.53 0.434 1.548 0.373 ;
        RECT 1.276 0.434 1.294 0.373 ;
        RECT 0.85 0.765 0.954 0.783 ;
        RECT 0.936 0.567 0.954 0.783 ;
        RECT 0.774 0.567 0.792 0.659 ;
        RECT 0.774 0.567 0.954 0.585 ;
        RECT 0.688 0.764 0.738 0.782 ;
        RECT 0.72 0.567 0.738 0.782 ;
        RECT 0.72 0.693 0.9 0.711 ;
        RECT 0.882 0.657 0.9 0.711 ;
        RECT 0.828 0.657 0.846 0.711 ;
        RECT 0.634 0.567 0.738 0.585 ;
        RECT 0.576 0.765 0.63 0.783 ;
        RECT 0.612 0.621 0.63 0.783 ;
        RECT 0.496 0.621 0.63 0.639 ;
        RECT 0.585 0.585 0.603 0.639 ;
        RECT 0.364 0.765 0.468 0.783 ;
        RECT 0.45 0.567 0.468 0.783 ;
        RECT 0.45 0.662 0.576 0.68 ;
        RECT 0.418 0.567 0.468 0.585 ;
        RECT 0.315 0.666 0.333 0.743 ;
        RECT 0.315 0.666 0.367 0.684 ;
        RECT 0.148 0.765 0.198 0.783 ;
        RECT 0.18 0.567 0.198 0.783 ;
        RECT 0.148 0.567 0.198 0.585 ;
        RECT 0.009 0.765 0.068 0.783 ;
        RECT 0.009 0.567 0.027 0.783 ;
        RECT 0.009 0.684 0.047 0.702 ;
        RECT 0.009 0.567 0.068 0.585 ;
        RECT 0.99 0.63 1.008 0.707 ;
        RECT 0.666 0.641 0.684 0.707 ;
        RECT 0.504 0.705 0.522 0.743 ;
        RECT 0.396 0.646 0.414 0.707 ;
        RECT 0.142 0.646 0.16 0.707 ;
        RECT 1.984 0.765 2.088 0.783 ;
        RECT 2.07 0.567 2.088 0.783 ;
        RECT 1.908 0.567 1.926 0.659 ;
        RECT 1.908 0.567 2.088 0.585 ;
        RECT 1.822 0.764 1.872 0.782 ;
        RECT 1.854 0.567 1.872 0.782 ;
        RECT 1.854 0.693 2.034 0.711 ;
        RECT 2.016 0.657 2.034 0.711 ;
        RECT 1.962 0.657 1.98 0.711 ;
        RECT 1.768 0.567 1.872 0.585 ;
        RECT 1.71 0.765 1.764 0.783 ;
        RECT 1.746 0.621 1.764 0.783 ;
        RECT 1.63 0.621 1.764 0.639 ;
        RECT 1.719 0.585 1.737 0.639 ;
        RECT 1.498 0.765 1.602 0.783 ;
        RECT 1.584 0.567 1.602 0.783 ;
        RECT 1.584 0.662 1.71 0.68 ;
        RECT 1.552 0.567 1.602 0.585 ;
        RECT 1.449 0.666 1.467 0.743 ;
        RECT 1.449 0.666 1.501 0.684 ;
        RECT 1.282 0.765 1.332 0.783 ;
        RECT 1.314 0.567 1.332 0.783 ;
        RECT 1.282 0.567 1.332 0.585 ;
        RECT 1.143 0.765 1.202 0.783 ;
        RECT 1.143 0.567 1.161 0.783 ;
        RECT 1.143 0.684 1.181 0.702 ;
        RECT 1.143 0.567 1.202 0.585 ;
        RECT 2.124 0.63 2.142 0.707 ;
        RECT 1.8 0.641 1.818 0.707 ;
        RECT 1.638 0.705 1.656 0.743 ;
        RECT 1.53 0.646 1.548 0.707 ;
        RECT 1.276 0.646 1.294 0.707 ;
        RECT 0.85 0.855 0.954 0.837 ;
        RECT 0.936 1.053 0.954 0.837 ;
        RECT 0.774 1.053 0.792 0.961 ;
        RECT 0.774 1.053 0.954 1.035 ;
        RECT 0.688 0.856 0.738 0.838 ;
        RECT 0.72 1.053 0.738 0.838 ;
        RECT 0.72 0.927 0.9 0.909 ;
        RECT 0.882 0.963 0.9 0.909 ;
        RECT 0.828 0.963 0.846 0.909 ;
        RECT 0.634 1.053 0.738 1.035 ;
        RECT 0.576 0.855 0.63 0.837 ;
        RECT 0.612 0.999 0.63 0.837 ;
        RECT 0.496 0.999 0.63 0.981 ;
        RECT 0.585 1.035 0.603 0.981 ;
        RECT 0.364 0.855 0.468 0.837 ;
        RECT 0.45 1.053 0.468 0.837 ;
        RECT 0.45 0.958 0.576 0.94 ;
        RECT 0.418 1.053 0.468 1.035 ;
        RECT 0.315 0.954 0.333 0.877 ;
        RECT 0.315 0.954 0.367 0.936 ;
        RECT 0.148 0.855 0.198 0.837 ;
        RECT 0.18 1.053 0.198 0.837 ;
        RECT 0.148 1.053 0.198 1.035 ;
        RECT 0.009 0.855 0.068 0.837 ;
        RECT 0.009 1.053 0.027 0.837 ;
        RECT 0.009 0.936 0.047 0.918 ;
        RECT 0.009 1.053 0.068 1.035 ;
        RECT 0.99 0.99 1.008 0.913 ;
        RECT 0.666 0.979 0.684 0.913 ;
        RECT 0.504 0.915 0.522 0.877 ;
        RECT 0.396 0.974 0.414 0.913 ;
        RECT 0.142 0.974 0.16 0.913 ;
        RECT 1.984 0.855 2.088 0.837 ;
        RECT 2.07 1.053 2.088 0.837 ;
        RECT 1.908 1.053 1.926 0.961 ;
        RECT 1.908 1.053 2.088 1.035 ;
        RECT 1.822 0.856 1.872 0.838 ;
        RECT 1.854 1.053 1.872 0.838 ;
        RECT 1.854 0.927 2.034 0.909 ;
        RECT 2.016 0.963 2.034 0.909 ;
        RECT 1.962 0.963 1.98 0.909 ;
        RECT 1.768 1.053 1.872 1.035 ;
        RECT 1.71 0.855 1.764 0.837 ;
        RECT 1.746 0.999 1.764 0.837 ;
        RECT 1.63 0.999 1.764 0.981 ;
        RECT 1.719 1.035 1.737 0.981 ;
        RECT 1.498 0.855 1.602 0.837 ;
        RECT 1.584 1.053 1.602 0.837 ;
        RECT 1.584 0.958 1.71 0.94 ;
        RECT 1.552 1.053 1.602 1.035 ;
        RECT 1.449 0.954 1.467 0.877 ;
        RECT 1.449 0.954 1.501 0.936 ;
        RECT 1.282 0.855 1.332 0.837 ;
        RECT 1.314 1.053 1.332 0.837 ;
        RECT 1.282 1.053 1.332 1.035 ;
        RECT 1.143 0.855 1.202 0.837 ;
        RECT 1.143 1.053 1.161 0.837 ;
        RECT 1.143 0.936 1.181 0.918 ;
        RECT 1.143 1.053 1.202 1.035 ;
        RECT 2.124 0.99 2.142 0.913 ;
        RECT 1.8 0.979 1.818 0.913 ;
        RECT 1.638 0.915 1.656 0.877 ;
        RECT 1.53 0.974 1.548 0.913 ;
        RECT 1.276 0.974 1.294 0.913 ;
        RECT 0.85 1.305 0.954 1.323 ;
        RECT 0.936 1.107 0.954 1.323 ;
        RECT 0.774 1.107 0.792 1.199 ;
        RECT 0.774 1.107 0.954 1.125 ;
        RECT 0.688 1.304 0.738 1.322 ;
        RECT 0.72 1.107 0.738 1.322 ;
        RECT 0.72 1.233 0.9 1.251 ;
        RECT 0.882 1.197 0.9 1.251 ;
        RECT 0.828 1.197 0.846 1.251 ;
        RECT 0.634 1.107 0.738 1.125 ;
        RECT 0.576 1.305 0.63 1.323 ;
        RECT 0.612 1.161 0.63 1.323 ;
        RECT 0.496 1.161 0.63 1.179 ;
        RECT 0.585 1.125 0.603 1.179 ;
        RECT 0.364 1.305 0.468 1.323 ;
        RECT 0.45 1.107 0.468 1.323 ;
        RECT 0.45 1.202 0.576 1.22 ;
        RECT 0.418 1.107 0.468 1.125 ;
        RECT 0.315 1.206 0.333 1.283 ;
        RECT 0.315 1.206 0.367 1.224 ;
        RECT 0.148 1.305 0.198 1.323 ;
        RECT 0.18 1.107 0.198 1.323 ;
        RECT 0.148 1.107 0.198 1.125 ;
        RECT 0.009 1.305 0.068 1.323 ;
        RECT 0.009 1.107 0.027 1.323 ;
        RECT 0.009 1.224 0.047 1.242 ;
        RECT 0.009 1.107 0.068 1.125 ;
        RECT 0.99 1.17 1.008 1.247 ;
        RECT 0.666 1.181 0.684 1.247 ;
        RECT 0.504 1.245 0.522 1.283 ;
        RECT 0.396 1.186 0.414 1.247 ;
        RECT 0.142 1.186 0.16 1.247 ;
        RECT 1.984 1.305 2.088 1.323 ;
        RECT 2.07 1.107 2.088 1.323 ;
        RECT 1.908 1.107 1.926 1.199 ;
        RECT 1.908 1.107 2.088 1.125 ;
        RECT 1.822 1.304 1.872 1.322 ;
        RECT 1.854 1.107 1.872 1.322 ;
        RECT 1.854 1.233 2.034 1.251 ;
        RECT 2.016 1.197 2.034 1.251 ;
        RECT 1.962 1.197 1.98 1.251 ;
        RECT 1.768 1.107 1.872 1.125 ;
        RECT 1.71 1.305 1.764 1.323 ;
        RECT 1.746 1.161 1.764 1.323 ;
        RECT 1.63 1.161 1.764 1.179 ;
        RECT 1.719 1.125 1.737 1.179 ;
        RECT 1.498 1.305 1.602 1.323 ;
        RECT 1.584 1.107 1.602 1.323 ;
        RECT 1.584 1.202 1.71 1.22 ;
        RECT 1.552 1.107 1.602 1.125 ;
        RECT 1.449 1.206 1.467 1.283 ;
        RECT 1.449 1.206 1.501 1.224 ;
        RECT 1.282 1.305 1.332 1.323 ;
        RECT 1.314 1.107 1.332 1.323 ;
        RECT 1.282 1.107 1.332 1.125 ;
        RECT 1.143 1.305 1.202 1.323 ;
        RECT 1.143 1.107 1.161 1.323 ;
        RECT 1.143 1.224 1.181 1.242 ;
        RECT 1.143 1.107 1.202 1.125 ;
        RECT 2.124 1.17 2.142 1.247 ;
        RECT 1.8 1.181 1.818 1.247 ;
        RECT 1.638 1.245 1.656 1.283 ;
        RECT 1.53 1.186 1.548 1.247 ;
        RECT 1.276 1.186 1.294 1.247 ;
        RECT 0.85 1.395 0.954 1.377 ;
        RECT 0.936 1.593 0.954 1.377 ;
        RECT 0.774 1.593 0.792 1.501 ;
        RECT 0.774 1.593 0.954 1.575 ;
        RECT 0.688 1.396 0.738 1.378 ;
        RECT 0.72 1.593 0.738 1.378 ;
        RECT 0.72 1.467 0.9 1.449 ;
        RECT 0.882 1.503 0.9 1.449 ;
        RECT 0.828 1.503 0.846 1.449 ;
        RECT 0.634 1.593 0.738 1.575 ;
        RECT 0.576 1.395 0.63 1.377 ;
        RECT 0.612 1.539 0.63 1.377 ;
        RECT 0.496 1.539 0.63 1.521 ;
        RECT 0.585 1.575 0.603 1.521 ;
        RECT 0.364 1.395 0.468 1.377 ;
        RECT 0.45 1.593 0.468 1.377 ;
        RECT 0.45 1.498 0.576 1.48 ;
        RECT 0.418 1.593 0.468 1.575 ;
        RECT 0.315 1.494 0.333 1.417 ;
        RECT 0.315 1.494 0.367 1.476 ;
        RECT 0.148 1.395 0.198 1.377 ;
        RECT 0.18 1.593 0.198 1.377 ;
        RECT 0.148 1.593 0.198 1.575 ;
        RECT 0.009 1.395 0.068 1.377 ;
        RECT 0.009 1.593 0.027 1.377 ;
        RECT 0.009 1.476 0.047 1.458 ;
        RECT 0.009 1.593 0.068 1.575 ;
        RECT 0.99 1.53 1.008 1.453 ;
        RECT 0.666 1.519 0.684 1.453 ;
        RECT 0.504 1.455 0.522 1.417 ;
        RECT 0.396 1.514 0.414 1.453 ;
        RECT 0.142 1.514 0.16 1.453 ;
        RECT 1.984 1.395 2.088 1.377 ;
        RECT 2.07 1.593 2.088 1.377 ;
        RECT 1.908 1.593 1.926 1.501 ;
        RECT 1.908 1.593 2.088 1.575 ;
        RECT 1.822 1.396 1.872 1.378 ;
        RECT 1.854 1.593 1.872 1.378 ;
        RECT 1.854 1.467 2.034 1.449 ;
        RECT 2.016 1.503 2.034 1.449 ;
        RECT 1.962 1.503 1.98 1.449 ;
        RECT 1.768 1.593 1.872 1.575 ;
        RECT 1.71 1.395 1.764 1.377 ;
        RECT 1.746 1.539 1.764 1.377 ;
        RECT 1.63 1.539 1.764 1.521 ;
        RECT 1.719 1.575 1.737 1.521 ;
        RECT 1.498 1.395 1.602 1.377 ;
        RECT 1.584 1.593 1.602 1.377 ;
        RECT 1.584 1.498 1.71 1.48 ;
        RECT 1.552 1.593 1.602 1.575 ;
        RECT 1.449 1.494 1.467 1.417 ;
        RECT 1.449 1.494 1.501 1.476 ;
        RECT 1.282 1.395 1.332 1.377 ;
        RECT 1.314 1.593 1.332 1.377 ;
        RECT 1.282 1.593 1.332 1.575 ;
        RECT 1.143 1.395 1.202 1.377 ;
        RECT 1.143 1.593 1.161 1.377 ;
        RECT 1.143 1.476 1.181 1.458 ;
        RECT 1.143 1.593 1.202 1.575 ;
        RECT 2.124 1.53 2.142 1.453 ;
        RECT 1.8 1.519 1.818 1.453 ;
        RECT 1.638 1.455 1.656 1.417 ;
        RECT 1.53 1.514 1.548 1.453 ;
        RECT 1.276 1.514 1.294 1.453 ;
        RECT 0.85 1.845 0.954 1.863 ;
        RECT 0.936 1.647 0.954 1.863 ;
        RECT 0.774 1.647 0.792 1.739 ;
        RECT 0.774 1.647 0.954 1.665 ;
        RECT 0.688 1.844 0.738 1.862 ;
        RECT 0.72 1.647 0.738 1.862 ;
        RECT 0.72 1.773 0.9 1.791 ;
        RECT 0.882 1.737 0.9 1.791 ;
        RECT 0.828 1.737 0.846 1.791 ;
        RECT 0.634 1.647 0.738 1.665 ;
        RECT 0.576 1.845 0.63 1.863 ;
        RECT 0.612 1.701 0.63 1.863 ;
        RECT 0.496 1.701 0.63 1.719 ;
        RECT 0.585 1.665 0.603 1.719 ;
        RECT 0.364 1.845 0.468 1.863 ;
        RECT 0.45 1.647 0.468 1.863 ;
        RECT 0.45 1.742 0.576 1.76 ;
        RECT 0.418 1.647 0.468 1.665 ;
        RECT 0.315 1.746 0.333 1.823 ;
        RECT 0.315 1.746 0.367 1.764 ;
        RECT 0.148 1.845 0.198 1.863 ;
        RECT 0.18 1.647 0.198 1.863 ;
        RECT 0.148 1.647 0.198 1.665 ;
        RECT 0.009 1.845 0.068 1.863 ;
        RECT 0.009 1.647 0.027 1.863 ;
        RECT 0.009 1.764 0.047 1.782 ;
        RECT 0.009 1.647 0.068 1.665 ;
        RECT 0.99 1.71 1.008 1.787 ;
        RECT 0.666 1.721 0.684 1.787 ;
        RECT 0.504 1.785 0.522 1.823 ;
        RECT 0.396 1.726 0.414 1.787 ;
        RECT 0.142 1.726 0.16 1.787 ;
        RECT 1.984 1.845 2.088 1.863 ;
        RECT 2.07 1.647 2.088 1.863 ;
        RECT 1.908 1.647 1.926 1.739 ;
        RECT 1.908 1.647 2.088 1.665 ;
        RECT 1.822 1.844 1.872 1.862 ;
        RECT 1.854 1.647 1.872 1.862 ;
        RECT 1.854 1.773 2.034 1.791 ;
        RECT 2.016 1.737 2.034 1.791 ;
        RECT 1.962 1.737 1.98 1.791 ;
        RECT 1.768 1.647 1.872 1.665 ;
        RECT 1.71 1.845 1.764 1.863 ;
        RECT 1.746 1.701 1.764 1.863 ;
        RECT 1.63 1.701 1.764 1.719 ;
        RECT 1.719 1.665 1.737 1.719 ;
        RECT 1.498 1.845 1.602 1.863 ;
        RECT 1.584 1.647 1.602 1.863 ;
        RECT 1.584 1.742 1.71 1.76 ;
        RECT 1.552 1.647 1.602 1.665 ;
        RECT 1.449 1.746 1.467 1.823 ;
        RECT 1.449 1.746 1.501 1.764 ;
        RECT 1.282 1.845 1.332 1.863 ;
        RECT 1.314 1.647 1.332 1.863 ;
        RECT 1.282 1.647 1.332 1.665 ;
        RECT 1.143 1.845 1.202 1.863 ;
        RECT 1.143 1.647 1.161 1.863 ;
        RECT 1.143 1.764 1.181 1.782 ;
        RECT 1.143 1.647 1.202 1.665 ;
        RECT 2.124 1.71 2.142 1.787 ;
        RECT 1.8 1.721 1.818 1.787 ;
        RECT 1.638 1.785 1.656 1.823 ;
        RECT 1.53 1.726 1.548 1.787 ;
        RECT 1.276 1.726 1.294 1.787 ;
        RECT 0.85 1.935 0.954 1.917 ;
        RECT 0.936 2.133 0.954 1.917 ;
        RECT 0.774 2.133 0.792 2.041 ;
        RECT 0.774 2.133 0.954 2.115 ;
        RECT 0.688 1.936 0.738 1.918 ;
        RECT 0.72 2.133 0.738 1.918 ;
        RECT 0.72 2.007 0.9 1.989 ;
        RECT 0.882 2.043 0.9 1.989 ;
        RECT 0.828 2.043 0.846 1.989 ;
        RECT 0.634 2.133 0.738 2.115 ;
        RECT 0.576 1.935 0.63 1.917 ;
        RECT 0.612 2.079 0.63 1.917 ;
        RECT 0.496 2.079 0.63 2.061 ;
        RECT 0.585 2.115 0.603 2.061 ;
        RECT 0.364 1.935 0.468 1.917 ;
        RECT 0.45 2.133 0.468 1.917 ;
        RECT 0.45 2.038 0.576 2.02 ;
        RECT 0.418 2.133 0.468 2.115 ;
        RECT 0.315 2.034 0.333 1.957 ;
        RECT 0.315 2.034 0.367 2.016 ;
        RECT 0.148 1.935 0.198 1.917 ;
        RECT 0.18 2.133 0.198 1.917 ;
        RECT 0.148 2.133 0.198 2.115 ;
        RECT 0.009 1.935 0.068 1.917 ;
        RECT 0.009 2.133 0.027 1.917 ;
        RECT 0.009 2.016 0.047 1.998 ;
        RECT 0.009 2.133 0.068 2.115 ;
        RECT 0.99 2.07 1.008 1.993 ;
        RECT 0.666 2.059 0.684 1.993 ;
        RECT 0.504 1.995 0.522 1.957 ;
        RECT 0.396 2.054 0.414 1.993 ;
        RECT 0.142 2.054 0.16 1.993 ;
        RECT 1.984 1.935 2.088 1.917 ;
        RECT 2.07 2.133 2.088 1.917 ;
        RECT 1.908 2.133 1.926 2.041 ;
        RECT 1.908 2.133 2.088 2.115 ;
        RECT 1.822 1.936 1.872 1.918 ;
        RECT 1.854 2.133 1.872 1.918 ;
        RECT 1.854 2.007 2.034 1.989 ;
        RECT 2.016 2.043 2.034 1.989 ;
        RECT 1.962 2.043 1.98 1.989 ;
        RECT 1.768 2.133 1.872 2.115 ;
        RECT 1.71 1.935 1.764 1.917 ;
        RECT 1.746 2.079 1.764 1.917 ;
        RECT 1.63 2.079 1.764 2.061 ;
        RECT 1.719 2.115 1.737 2.061 ;
        RECT 1.498 1.935 1.602 1.917 ;
        RECT 1.584 2.133 1.602 1.917 ;
        RECT 1.584 2.038 1.71 2.02 ;
        RECT 1.552 2.133 1.602 2.115 ;
        RECT 1.449 2.034 1.467 1.957 ;
        RECT 1.449 2.034 1.501 2.016 ;
        RECT 1.282 1.935 1.332 1.917 ;
        RECT 1.314 2.133 1.332 1.917 ;
        RECT 1.282 2.133 1.332 2.115 ;
        RECT 1.143 1.935 1.202 1.917 ;
        RECT 1.143 2.133 1.161 1.917 ;
        RECT 1.143 2.016 1.181 1.998 ;
        RECT 1.143 2.133 1.202 2.115 ;
        RECT 2.124 2.07 2.142 1.993 ;
        RECT 1.8 2.059 1.818 1.993 ;
        RECT 1.638 1.995 1.656 1.957 ;
        RECT 1.53 2.054 1.548 1.993 ;
        RECT 1.276 2.054 1.294 1.993 ;
      LAYER M2 ;
        RECT 0.877 0.144 1.013 0.162 ;
        RECT 0.019 0.144 0.689 0.162 ;
        RECT 0.175 0.18 0.527 0.198 ;
        RECT 2.011 0.144 2.147 0.162 ;
        RECT 1.153 0.144 1.823 0.162 ;
        RECT 1.309 0.18 1.661 0.198 ;
        RECT 0.877 0.396 1.013 0.378 ;
        RECT 0.019 0.396 0.689 0.378 ;
        RECT 0.175 0.36 0.527 0.342 ;
        RECT 2.011 0.396 2.147 0.378 ;
        RECT 1.153 0.396 1.823 0.378 ;
        RECT 1.309 0.36 1.661 0.342 ;
        RECT 0.877 0.684 1.013 0.702 ;
        RECT 0.019 0.684 0.689 0.702 ;
        RECT 0.175 0.72 0.527 0.738 ;
        RECT 2.011 0.684 2.147 0.702 ;
        RECT 1.153 0.684 1.823 0.702 ;
        RECT 1.309 0.72 1.661 0.738 ;
        RECT 0.877 0.936 1.013 0.918 ;
        RECT 0.019 0.936 0.689 0.918 ;
        RECT 0.175 0.9 0.527 0.882 ;
        RECT 2.011 0.936 2.147 0.918 ;
        RECT 1.153 0.936 1.823 0.918 ;
        RECT 1.309 0.9 1.661 0.882 ;
        RECT 0.877 1.224 1.013 1.242 ;
        RECT 0.019 1.224 0.689 1.242 ;
        RECT 0.175 1.26 0.527 1.278 ;
        RECT 2.011 1.224 2.147 1.242 ;
        RECT 1.153 1.224 1.823 1.242 ;
        RECT 1.309 1.26 1.661 1.278 ;
        RECT 0.877 1.476 1.013 1.458 ;
        RECT 0.019 1.476 0.689 1.458 ;
        RECT 0.175 1.44 0.527 1.422 ;
        RECT 2.011 1.476 2.147 1.458 ;
        RECT 1.153 1.476 1.823 1.458 ;
        RECT 1.309 1.44 1.661 1.422 ;
        RECT 0.877 1.764 1.013 1.782 ;
        RECT 0.019 1.764 0.689 1.782 ;
        RECT 0.175 1.8 0.527 1.818 ;
        RECT 2.011 1.764 2.147 1.782 ;
        RECT 1.153 1.764 1.823 1.782 ;
        RECT 1.309 1.8 1.661 1.818 ;
        RECT 0.877 2.016 1.013 1.998 ;
        RECT 0.019 2.016 0.689 1.998 ;
        RECT 0.175 1.98 0.527 1.962 ;
        RECT 2.011 2.016 2.147 1.998 ;
        RECT 1.153 2.016 1.823 1.998 ;
        RECT 1.309 1.98 1.661 1.962 ;
      LAYER V1 ;
        RECT 0.99 0.144 1.008 0.162 ;
        RECT 0.882 0.144 0.9 0.162 ;
        RECT 0.666 0.144 0.684 0.162 ;
        RECT 0.504 0.18 0.522 0.198 ;
        RECT 0.396 0.144 0.414 0.162 ;
        RECT 0.315 0.18 0.333 0.198 ;
        RECT 0.18 0.18 0.198 0.198 ;
        RECT 0.142 0.144 0.16 0.162 ;
        RECT 0.024 0.144 0.042 0.162 ;
        RECT 2.124 0.144 2.142 0.162 ;
        RECT 2.016 0.144 2.034 0.162 ;
        RECT 1.8 0.144 1.818 0.162 ;
        RECT 1.638 0.18 1.656 0.198 ;
        RECT 1.53 0.144 1.548 0.162 ;
        RECT 1.449 0.18 1.467 0.198 ;
        RECT 1.314 0.18 1.332 0.198 ;
        RECT 1.276 0.144 1.294 0.162 ;
        RECT 1.158 0.144 1.176 0.162 ;
        RECT 0.99 0.396 1.008 0.378 ;
        RECT 0.882 0.396 0.9 0.378 ;
        RECT 0.666 0.396 0.684 0.378 ;
        RECT 0.504 0.36 0.522 0.342 ;
        RECT 0.396 0.396 0.414 0.378 ;
        RECT 0.315 0.36 0.333 0.342 ;
        RECT 0.18 0.36 0.198 0.342 ;
        RECT 0.142 0.396 0.16 0.378 ;
        RECT 0.024 0.396 0.042 0.378 ;
        RECT 2.124 0.396 2.142 0.378 ;
        RECT 2.016 0.396 2.034 0.378 ;
        RECT 1.8 0.396 1.818 0.378 ;
        RECT 1.638 0.36 1.656 0.342 ;
        RECT 1.53 0.396 1.548 0.378 ;
        RECT 1.449 0.36 1.467 0.342 ;
        RECT 1.314 0.36 1.332 0.342 ;
        RECT 1.276 0.396 1.294 0.378 ;
        RECT 1.158 0.396 1.176 0.378 ;
        RECT 0.99 0.684 1.008 0.702 ;
        RECT 0.882 0.684 0.9 0.702 ;
        RECT 0.666 0.684 0.684 0.702 ;
        RECT 0.504 0.72 0.522 0.738 ;
        RECT 0.396 0.684 0.414 0.702 ;
        RECT 0.315 0.72 0.333 0.738 ;
        RECT 0.18 0.72 0.198 0.738 ;
        RECT 0.142 0.684 0.16 0.702 ;
        RECT 0.024 0.684 0.042 0.702 ;
        RECT 2.124 0.684 2.142 0.702 ;
        RECT 2.016 0.684 2.034 0.702 ;
        RECT 1.8 0.684 1.818 0.702 ;
        RECT 1.638 0.72 1.656 0.738 ;
        RECT 1.53 0.684 1.548 0.702 ;
        RECT 1.449 0.72 1.467 0.738 ;
        RECT 1.314 0.72 1.332 0.738 ;
        RECT 1.276 0.684 1.294 0.702 ;
        RECT 1.158 0.684 1.176 0.702 ;
        RECT 0.99 0.936 1.008 0.918 ;
        RECT 0.882 0.936 0.9 0.918 ;
        RECT 0.666 0.936 0.684 0.918 ;
        RECT 0.504 0.9 0.522 0.882 ;
        RECT 0.396 0.936 0.414 0.918 ;
        RECT 0.315 0.9 0.333 0.882 ;
        RECT 0.18 0.9 0.198 0.882 ;
        RECT 0.142 0.936 0.16 0.918 ;
        RECT 0.024 0.936 0.042 0.918 ;
        RECT 2.124 0.936 2.142 0.918 ;
        RECT 2.016 0.936 2.034 0.918 ;
        RECT 1.8 0.936 1.818 0.918 ;
        RECT 1.638 0.9 1.656 0.882 ;
        RECT 1.53 0.936 1.548 0.918 ;
        RECT 1.449 0.9 1.467 0.882 ;
        RECT 1.314 0.9 1.332 0.882 ;
        RECT 1.276 0.936 1.294 0.918 ;
        RECT 1.158 0.936 1.176 0.918 ;
        RECT 0.99 1.224 1.008 1.242 ;
        RECT 0.882 1.224 0.9 1.242 ;
        RECT 0.666 1.224 0.684 1.242 ;
        RECT 0.504 1.26 0.522 1.278 ;
        RECT 0.396 1.224 0.414 1.242 ;
        RECT 0.315 1.26 0.333 1.278 ;
        RECT 0.18 1.26 0.198 1.278 ;
        RECT 0.142 1.224 0.16 1.242 ;
        RECT 0.024 1.224 0.042 1.242 ;
        RECT 2.124 1.224 2.142 1.242 ;
        RECT 2.016 1.224 2.034 1.242 ;
        RECT 1.8 1.224 1.818 1.242 ;
        RECT 1.638 1.26 1.656 1.278 ;
        RECT 1.53 1.224 1.548 1.242 ;
        RECT 1.449 1.26 1.467 1.278 ;
        RECT 1.314 1.26 1.332 1.278 ;
        RECT 1.276 1.224 1.294 1.242 ;
        RECT 1.158 1.224 1.176 1.242 ;
        RECT 0.99 1.476 1.008 1.458 ;
        RECT 0.882 1.476 0.9 1.458 ;
        RECT 0.666 1.476 0.684 1.458 ;
        RECT 0.504 1.44 0.522 1.422 ;
        RECT 0.396 1.476 0.414 1.458 ;
        RECT 0.315 1.44 0.333 1.422 ;
        RECT 0.18 1.44 0.198 1.422 ;
        RECT 0.142 1.476 0.16 1.458 ;
        RECT 0.024 1.476 0.042 1.458 ;
        RECT 2.124 1.476 2.142 1.458 ;
        RECT 2.016 1.476 2.034 1.458 ;
        RECT 1.8 1.476 1.818 1.458 ;
        RECT 1.638 1.44 1.656 1.422 ;
        RECT 1.53 1.476 1.548 1.458 ;
        RECT 1.449 1.44 1.467 1.422 ;
        RECT 1.314 1.44 1.332 1.422 ;
        RECT 1.276 1.476 1.294 1.458 ;
        RECT 1.158 1.476 1.176 1.458 ;
        RECT 0.99 1.764 1.008 1.782 ;
        RECT 0.882 1.764 0.9 1.782 ;
        RECT 0.666 1.764 0.684 1.782 ;
        RECT 0.504 1.8 0.522 1.818 ;
        RECT 0.396 1.764 0.414 1.782 ;
        RECT 0.315 1.8 0.333 1.818 ;
        RECT 0.18 1.8 0.198 1.818 ;
        RECT 0.142 1.764 0.16 1.782 ;
        RECT 0.024 1.764 0.042 1.782 ;
        RECT 2.124 1.764 2.142 1.782 ;
        RECT 2.016 1.764 2.034 1.782 ;
        RECT 1.8 1.764 1.818 1.782 ;
        RECT 1.638 1.8 1.656 1.818 ;
        RECT 1.53 1.764 1.548 1.782 ;
        RECT 1.449 1.8 1.467 1.818 ;
        RECT 1.314 1.8 1.332 1.818 ;
        RECT 1.276 1.764 1.294 1.782 ;
        RECT 1.158 1.764 1.176 1.782 ;
        RECT 0.99 2.016 1.008 1.998 ;
        RECT 0.882 2.016 0.9 1.998 ;
        RECT 0.666 2.016 0.684 1.998 ;
        RECT 0.504 1.98 0.522 1.962 ;
        RECT 0.396 2.016 0.414 1.998 ;
        RECT 0.315 1.98 0.333 1.962 ;
        RECT 0.18 1.98 0.198 1.962 ;
        RECT 0.142 2.016 0.16 1.998 ;
        RECT 0.024 2.016 0.042 1.998 ;
        RECT 2.124 2.016 2.142 1.998 ;
        RECT 2.016 2.016 2.034 1.998 ;
        RECT 1.8 2.016 1.818 1.998 ;
        RECT 1.638 1.98 1.656 1.962 ;
        RECT 1.53 2.016 1.548 1.998 ;
        RECT 1.449 1.98 1.467 1.962 ;
        RECT 1.314 1.98 1.332 1.962 ;
        RECT 1.276 2.016 1.294 1.998 ;
        RECT 1.158 2.016 1.176 1.998 ;
    END
END DFFHQNV8H2Xx2_ASAP7_75t_SL

END LIBRARY
