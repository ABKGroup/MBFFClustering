VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_1024x39
  FOREIGN fakeram7_1024x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 20.330 BY 67.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.768 0.024 0.792 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.112 0.024 2.136 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.784 0.024 2.808 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.456 0.024 3.480 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.800 0.024 4.824 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.144 0.024 6.168 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.816 0.024 6.840 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.160 0.024 8.184 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.832 0.024 8.856 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.504 0.024 9.528 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.176 0.024 10.200 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.848 0.024 10.872 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.520 0.024 11.544 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.192 0.024 12.216 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.864 0.024 12.888 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.536 0.024 13.560 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.208 0.024 14.232 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.880 0.024 14.904 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.552 0.024 15.576 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.224 0.024 16.248 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.896 0.024 16.920 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.568 0.024 17.592 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.240 0.024 18.264 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.912 0.024 18.936 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.584 0.024 19.608 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.256 0.024 20.280 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.928 0.024 20.952 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.600 0.024 21.624 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.272 0.024 22.296 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.944 0.024 22.968 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.616 0.024 23.640 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.288 0.024 24.312 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.960 0.024 24.984 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.632 0.024 25.656 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.072 0.024 27.096 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.744 0.024 27.768 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.416 0.024 28.440 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.088 0.024 29.112 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.760 0.024 29.784 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.432 0.024 30.456 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.104 0.024 31.128 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.776 0.024 31.800 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.448 0.024 32.472 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.120 0.024 33.144 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.792 0.024 33.816 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.464 0.024 34.488 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.136 0.024 35.160 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.808 0.024 35.832 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.480 0.024 36.504 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.152 0.024 37.176 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.824 0.024 37.848 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.496 0.024 38.520 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.168 0.024 39.192 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.840 0.024 39.864 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.512 0.024 40.536 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.184 0.024 41.208 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.856 0.024 41.880 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.528 0.024 42.552 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.200 0.024 43.224 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.872 0.024 43.896 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.544 0.024 44.568 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.216 0.024 45.240 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.888 0.024 45.912 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.560 0.024 46.584 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.232 0.024 47.256 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.904 0.024 47.928 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.576 0.024 48.600 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.248 0.024 49.272 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.920 0.024 49.944 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.592 0.024 50.616 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.264 0.024 51.288 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.936 0.024 51.960 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.608 0.024 52.632 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.048 0.024 54.072 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.720 0.024 54.744 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.392 0.024 55.416 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.064 0.024 56.088 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.736 0.024 56.760 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.408 0.024 57.432 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.080 0.024 58.104 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.752 0.024 58.776 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.424 0.024 59.448 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.096 0.024 60.120 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.536 0.024 61.560 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.208 0.024 62.232 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.880 0.024 62.904 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 20.234 0.144 ;
      RECT 0.096 1.584 20.234 1.680 ;
      RECT 0.096 3.120 20.234 3.216 ;
      RECT 0.096 4.656 20.234 4.752 ;
      RECT 0.096 6.192 20.234 6.288 ;
      RECT 0.096 7.728 20.234 7.824 ;
      RECT 0.096 9.264 20.234 9.360 ;
      RECT 0.096 10.800 20.234 10.896 ;
      RECT 0.096 12.336 20.234 12.432 ;
      RECT 0.096 13.872 20.234 13.968 ;
      RECT 0.096 15.408 20.234 15.504 ;
      RECT 0.096 16.944 20.234 17.040 ;
      RECT 0.096 18.480 20.234 18.576 ;
      RECT 0.096 20.016 20.234 20.112 ;
      RECT 0.096 21.552 20.234 21.648 ;
      RECT 0.096 23.088 20.234 23.184 ;
      RECT 0.096 24.624 20.234 24.720 ;
      RECT 0.096 26.160 20.234 26.256 ;
      RECT 0.096 27.696 20.234 27.792 ;
      RECT 0.096 29.232 20.234 29.328 ;
      RECT 0.096 30.768 20.234 30.864 ;
      RECT 0.096 32.304 20.234 32.400 ;
      RECT 0.096 33.840 20.234 33.936 ;
      RECT 0.096 35.376 20.234 35.472 ;
      RECT 0.096 36.912 20.234 37.008 ;
      RECT 0.096 38.448 20.234 38.544 ;
      RECT 0.096 39.984 20.234 40.080 ;
      RECT 0.096 41.520 20.234 41.616 ;
      RECT 0.096 43.056 20.234 43.152 ;
      RECT 0.096 44.592 20.234 44.688 ;
      RECT 0.096 46.128 20.234 46.224 ;
      RECT 0.096 47.664 20.234 47.760 ;
      RECT 0.096 49.200 20.234 49.296 ;
      RECT 0.096 50.736 20.234 50.832 ;
      RECT 0.096 52.272 20.234 52.368 ;
      RECT 0.096 53.808 20.234 53.904 ;
      RECT 0.096 55.344 20.234 55.440 ;
      RECT 0.096 56.880 20.234 56.976 ;
      RECT 0.096 58.416 20.234 58.512 ;
      RECT 0.096 59.952 20.234 60.048 ;
      RECT 0.096 61.488 20.234 61.584 ;
      RECT 0.096 63.024 20.234 63.120 ;
      RECT 0.096 64.560 20.234 64.656 ;
      RECT 0.096 66.096 20.234 66.192 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 20.234 0.912 ;
      RECT 0.096 2.352 20.234 2.448 ;
      RECT 0.096 3.888 20.234 3.984 ;
      RECT 0.096 5.424 20.234 5.520 ;
      RECT 0.096 6.960 20.234 7.056 ;
      RECT 0.096 8.496 20.234 8.592 ;
      RECT 0.096 10.032 20.234 10.128 ;
      RECT 0.096 11.568 20.234 11.664 ;
      RECT 0.096 13.104 20.234 13.200 ;
      RECT 0.096 14.640 20.234 14.736 ;
      RECT 0.096 16.176 20.234 16.272 ;
      RECT 0.096 17.712 20.234 17.808 ;
      RECT 0.096 19.248 20.234 19.344 ;
      RECT 0.096 20.784 20.234 20.880 ;
      RECT 0.096 22.320 20.234 22.416 ;
      RECT 0.096 23.856 20.234 23.952 ;
      RECT 0.096 25.392 20.234 25.488 ;
      RECT 0.096 26.928 20.234 27.024 ;
      RECT 0.096 28.464 20.234 28.560 ;
      RECT 0.096 30.000 20.234 30.096 ;
      RECT 0.096 31.536 20.234 31.632 ;
      RECT 0.096 33.072 20.234 33.168 ;
      RECT 0.096 34.608 20.234 34.704 ;
      RECT 0.096 36.144 20.234 36.240 ;
      RECT 0.096 37.680 20.234 37.776 ;
      RECT 0.096 39.216 20.234 39.312 ;
      RECT 0.096 40.752 20.234 40.848 ;
      RECT 0.096 42.288 20.234 42.384 ;
      RECT 0.096 43.824 20.234 43.920 ;
      RECT 0.096 45.360 20.234 45.456 ;
      RECT 0.096 46.896 20.234 46.992 ;
      RECT 0.096 48.432 20.234 48.528 ;
      RECT 0.096 49.968 20.234 50.064 ;
      RECT 0.096 51.504 20.234 51.600 ;
      RECT 0.096 53.040 20.234 53.136 ;
      RECT 0.096 54.576 20.234 54.672 ;
      RECT 0.096 56.112 20.234 56.208 ;
      RECT 0.096 57.648 20.234 57.744 ;
      RECT 0.096 59.184 20.234 59.280 ;
      RECT 0.096 60.720 20.234 60.816 ;
      RECT 0.096 62.256 20.234 62.352 ;
      RECT 0.096 63.792 20.234 63.888 ;
      RECT 0.096 65.328 20.234 65.424 ;
      RECT 0.096 66.864 20.234 66.960 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 20.330 67.200 ;
    LAYER M2 ;
    RECT 0 0 20.330 67.200 ;
    LAYER M3 ;
    RECT 0 0 20.330 67.200 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 67.200 ;
    RECT 20.234 0 20.330 67.200 ;
    RECT 0.096 0.000 20.234 0.048 ;
    RECT 0.096 0.144 20.234 0.816 ;
    RECT 0.096 0.912 20.234 1.584 ;
    RECT 0.096 1.680 20.234 2.352 ;
    RECT 0.096 2.448 20.234 3.120 ;
    RECT 0.096 3.216 20.234 3.888 ;
    RECT 0.096 3.984 20.234 4.656 ;
    RECT 0.096 4.752 20.234 5.424 ;
    RECT 0.096 5.520 20.234 6.192 ;
    RECT 0.096 6.288 20.234 6.960 ;
    RECT 0.096 7.056 20.234 7.728 ;
    RECT 0.096 7.824 20.234 8.496 ;
    RECT 0.096 8.592 20.234 9.264 ;
    RECT 0.096 9.360 20.234 10.032 ;
    RECT 0.096 10.128 20.234 10.800 ;
    RECT 0.096 10.896 20.234 11.568 ;
    RECT 0.096 11.664 20.234 12.336 ;
    RECT 0.096 12.432 20.234 13.104 ;
    RECT 0.096 13.200 20.234 13.872 ;
    RECT 0.096 13.968 20.234 14.640 ;
    RECT 0.096 14.736 20.234 15.408 ;
    RECT 0.096 15.504 20.234 16.176 ;
    RECT 0.096 16.272 20.234 16.944 ;
    RECT 0.096 17.040 20.234 17.712 ;
    RECT 0.096 17.808 20.234 18.480 ;
    RECT 0.096 18.576 20.234 19.248 ;
    RECT 0.096 19.344 20.234 20.016 ;
    RECT 0.096 20.112 20.234 20.784 ;
    RECT 0.096 20.880 20.234 21.552 ;
    RECT 0.096 21.648 20.234 22.320 ;
    RECT 0.096 22.416 20.234 23.088 ;
    RECT 0.096 23.184 20.234 23.856 ;
    RECT 0.096 23.952 20.234 24.624 ;
    RECT 0.096 24.720 20.234 25.392 ;
    RECT 0.096 25.488 20.234 26.160 ;
    RECT 0.096 26.256 20.234 26.928 ;
    RECT 0.096 27.024 20.234 27.696 ;
    RECT 0.096 27.792 20.234 28.464 ;
    RECT 0.096 28.560 20.234 29.232 ;
    RECT 0.096 29.328 20.234 30.000 ;
    RECT 0.096 30.096 20.234 30.768 ;
    RECT 0.096 30.864 20.234 31.536 ;
    RECT 0.096 31.632 20.234 32.304 ;
    RECT 0.096 32.400 20.234 33.072 ;
    RECT 0.096 33.168 20.234 33.840 ;
    RECT 0.096 33.936 20.234 34.608 ;
    RECT 0.096 34.704 20.234 35.376 ;
    RECT 0.096 35.472 20.234 36.144 ;
    RECT 0.096 36.240 20.234 36.912 ;
    RECT 0.096 37.008 20.234 37.680 ;
    RECT 0.096 37.776 20.234 38.448 ;
    RECT 0.096 38.544 20.234 39.216 ;
    RECT 0.096 39.312 20.234 39.984 ;
    RECT 0.096 40.080 20.234 40.752 ;
    RECT 0.096 40.848 20.234 41.520 ;
    RECT 0.096 41.616 20.234 42.288 ;
    RECT 0.096 42.384 20.234 43.056 ;
    RECT 0.096 43.152 20.234 43.824 ;
    RECT 0.096 43.920 20.234 44.592 ;
    RECT 0.096 44.688 20.234 45.360 ;
    RECT 0.096 45.456 20.234 46.128 ;
    RECT 0.096 46.224 20.234 46.896 ;
    RECT 0.096 46.992 20.234 47.664 ;
    RECT 0.096 47.760 20.234 48.432 ;
    RECT 0.096 48.528 20.234 49.200 ;
    RECT 0.096 49.296 20.234 49.968 ;
    RECT 0.096 50.064 20.234 50.736 ;
    RECT 0.096 50.832 20.234 51.504 ;
    RECT 0.096 51.600 20.234 52.272 ;
    RECT 0.096 52.368 20.234 53.040 ;
    RECT 0.096 53.136 20.234 53.808 ;
    RECT 0.096 53.904 20.234 54.576 ;
    RECT 0.096 54.672 20.234 55.344 ;
    RECT 0.096 55.440 20.234 56.112 ;
    RECT 0.096 56.208 20.234 56.880 ;
    RECT 0.096 56.976 20.234 57.648 ;
    RECT 0.096 57.744 20.234 58.416 ;
    RECT 0.096 58.512 20.234 59.184 ;
    RECT 0.096 59.280 20.234 59.952 ;
    RECT 0.096 60.048 20.234 60.720 ;
    RECT 0.096 60.816 20.234 61.488 ;
    RECT 0.096 61.584 20.234 62.256 ;
    RECT 0.096 62.352 20.234 63.024 ;
    RECT 0.096 63.120 20.234 63.792 ;
    RECT 0.096 63.888 20.234 64.560 ;
    RECT 0.096 64.656 20.234 65.328 ;
    RECT 0.096 65.424 20.234 66.096 ;
    RECT 0.096 66.192 20.234 66.864 ;
    RECT 0.096 66.960 20.234 67.200 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 0.768 ;
    RECT 0 0.792 0.024 1.440 ;
    RECT 0 1.464 0.024 2.112 ;
    RECT 0 2.136 0.024 2.784 ;
    RECT 0 2.808 0.024 3.456 ;
    RECT 0 3.480 0.024 4.128 ;
    RECT 0 4.152 0.024 4.800 ;
    RECT 0 4.824 0.024 5.472 ;
    RECT 0 5.496 0.024 6.144 ;
    RECT 0 6.168 0.024 6.816 ;
    RECT 0 6.840 0.024 7.488 ;
    RECT 0 7.512 0.024 8.160 ;
    RECT 0 8.184 0.024 8.832 ;
    RECT 0 8.856 0.024 9.504 ;
    RECT 0 9.528 0.024 10.176 ;
    RECT 0 10.200 0.024 10.848 ;
    RECT 0 10.872 0.024 11.520 ;
    RECT 0 11.544 0.024 12.192 ;
    RECT 0 12.216 0.024 12.864 ;
    RECT 0 12.888 0.024 13.536 ;
    RECT 0 13.560 0.024 14.208 ;
    RECT 0 14.232 0.024 14.880 ;
    RECT 0 14.904 0.024 15.552 ;
    RECT 0 15.576 0.024 16.224 ;
    RECT 0 16.248 0.024 16.896 ;
    RECT 0 16.920 0.024 17.568 ;
    RECT 0 17.592 0.024 18.240 ;
    RECT 0 18.264 0.024 18.912 ;
    RECT 0 18.936 0.024 19.584 ;
    RECT 0 19.608 0.024 20.256 ;
    RECT 0 20.280 0.024 20.928 ;
    RECT 0 20.952 0.024 21.600 ;
    RECT 0 21.624 0.024 22.272 ;
    RECT 0 22.296 0.024 22.944 ;
    RECT 0 22.968 0.024 23.616 ;
    RECT 0 23.640 0.024 24.288 ;
    RECT 0 24.312 0.024 24.960 ;
    RECT 0 24.984 0.024 25.632 ;
    RECT 0 25.656 0.024 27.072 ;
    RECT 0 27.096 0.024 27.744 ;
    RECT 0 27.768 0.024 28.416 ;
    RECT 0 28.440 0.024 29.088 ;
    RECT 0 29.112 0.024 29.760 ;
    RECT 0 29.784 0.024 30.432 ;
    RECT 0 30.456 0.024 31.104 ;
    RECT 0 31.128 0.024 31.776 ;
    RECT 0 31.800 0.024 32.448 ;
    RECT 0 32.472 0.024 33.120 ;
    RECT 0 33.144 0.024 33.792 ;
    RECT 0 33.816 0.024 34.464 ;
    RECT 0 34.488 0.024 35.136 ;
    RECT 0 35.160 0.024 35.808 ;
    RECT 0 35.832 0.024 36.480 ;
    RECT 0 36.504 0.024 37.152 ;
    RECT 0 37.176 0.024 37.824 ;
    RECT 0 37.848 0.024 38.496 ;
    RECT 0 38.520 0.024 39.168 ;
    RECT 0 39.192 0.024 39.840 ;
    RECT 0 39.864 0.024 40.512 ;
    RECT 0 40.536 0.024 41.184 ;
    RECT 0 41.208 0.024 41.856 ;
    RECT 0 41.880 0.024 42.528 ;
    RECT 0 42.552 0.024 43.200 ;
    RECT 0 43.224 0.024 43.872 ;
    RECT 0 43.896 0.024 44.544 ;
    RECT 0 44.568 0.024 45.216 ;
    RECT 0 45.240 0.024 45.888 ;
    RECT 0 45.912 0.024 46.560 ;
    RECT 0 46.584 0.024 47.232 ;
    RECT 0 47.256 0.024 47.904 ;
    RECT 0 47.928 0.024 48.576 ;
    RECT 0 48.600 0.024 49.248 ;
    RECT 0 49.272 0.024 49.920 ;
    RECT 0 49.944 0.024 50.592 ;
    RECT 0 50.616 0.024 51.264 ;
    RECT 0 51.288 0.024 51.936 ;
    RECT 0 51.960 0.024 52.608 ;
    RECT 0 52.632 0.024 54.048 ;
    RECT 0 54.072 0.024 54.720 ;
    RECT 0 54.744 0.024 55.392 ;
    RECT 0 55.416 0.024 56.064 ;
    RECT 0 56.088 0.024 56.736 ;
    RECT 0 56.760 0.024 57.408 ;
    RECT 0 57.432 0.024 58.080 ;
    RECT 0 58.104 0.024 58.752 ;
    RECT 0 58.776 0.024 59.424 ;
    RECT 0 59.448 0.024 60.096 ;
    RECT 0 60.120 0.024 60.768 ;
    RECT 0 60.792 0.024 61.440 ;
    RECT 0 61.464 0.024 62.112 ;
    RECT 0 62.136 0.024 62.784 ;
    RECT 0 62.808 0.024 63.456 ;
    RECT 0 63.480 0.024 64.128 ;
    RECT 0 64.152 0.024 64.800 ;
    RECT 0 64.824 0.024 65.472 ;
    RECT 0 65.496 0.024 66.144 ;
    RECT 0 66.168 0.024 66.816 ;
    RECT 0 66.840 0.024 67.488 ;
    RECT 0 67.512 0.024 68.160 ;
    RECT 0 68.184 0.024 68.832 ;
    RECT 0 68.856 0.024 69.504 ;
    RECT 0 69.528 0.024 70.176 ;
    RECT 0 70.200 0.024 70.848 ;
    RECT 0 70.872 0.024 71.520 ;
    RECT 0 71.544 0.024 72.192 ;
    RECT 0 72.216 0.024 72.864 ;
    RECT 0 72.888 0.024 73.536 ;
    RECT 0 73.560 0.024 74.208 ;
    RECT 0 74.232 0.024 74.880 ;
    RECT 0 74.904 0.024 75.552 ;
    RECT 0 75.576 0.024 76.224 ;
    RECT 0 76.248 0.024 76.896 ;
    RECT 0 76.920 0.024 77.568 ;
    RECT 0 77.592 0.024 78.240 ;
    RECT 0 78.264 0.024 78.912 ;
    RECT 0 78.936 0.024 79.584 ;
    RECT 0 79.608 0.024 81.024 ;
    RECT 0 81.048 0.024 81.696 ;
    RECT 0 81.720 0.024 82.368 ;
    RECT 0 82.392 0.024 83.040 ;
    RECT 0 83.064 0.024 83.712 ;
    RECT 0 83.736 0.024 84.384 ;
    RECT 0 84.408 0.024 85.056 ;
    RECT 0 85.080 0.024 85.728 ;
    RECT 0 85.752 0.024 86.400 ;
    RECT 0 86.424 0.024 87.072 ;
    RECT 0 87.096 0.024 88.512 ;
    RECT 0 88.536 0.024 89.184 ;
    RECT 0 89.208 0.024 89.856 ;
    RECT 0 89.880 0.024 67.200 ;
    LAYER OVERLAP ;
    RECT 0 0 20.330 67.200 ;
  END
END fakeram7_1024x39

END LIBRARY
