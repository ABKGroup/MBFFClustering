VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE asap7sc7p5t_R8
  CLASS CORE ;
  SIZE 0.054 BY 2.16 ;
  SYMMETRY Y ;
END asap7sc7p5t_R8

MACRO DFFHQNV8H2Xx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0.0 0.0 ;
  FOREIGN DFFHQNV8H2Xx1_ASAP7_75t_L 0.0 0.0 ;
  SIZE 2.16 BY 2.16 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_R8 ;
    PIN VDD
      USE POWER ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 0.261 1.08 0.279 ;
          RECT 1.08 0.261 2.16 0.279 ;
          RECT 0.0 0.801 1.08 0.819 ;
          RECT 1.08 0.801 2.16 0.819 ;
          RECT 0.0 1.341 1.08 1.359 ;
          RECT 1.08 1.341 2.16 1.359 ;
          RECT 0.0 1.881 1.08 1.899 ;
          RECT 1.08 1.881 2.16 1.899 ;
      END
    END VDD
    PIN VSS
      USE GROUND ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 -0.009 1.08 0.009 ;
          RECT 1.08 -0.009 2.16 0.009 ;
          RECT 0.0 0.549 1.08 0.531 ;
          RECT 1.08 0.549 2.16 0.531 ;
          RECT 0.0 1.089 1.08 1.071 ;
          RECT 1.08 1.089 2.16 1.071 ;
          RECT 0.0 1.629 1.08 1.611 ;
          RECT 1.08 1.629 2.16 1.611 ;
          RECT 0.0 2.169 1.08 2.151 ;
          RECT 1.08 2.169 2.16 2.151 ;
      END
    END VSS
    PIN CLK
      USE CLOCK ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.099 0.164 0.117 0.236 ;
          RECT 0.072 0.07 0.117 0.106 ;
          RECT 0.099 0.034 0.117 0.106 ;
          RECT 0.072 0.164 0.117 0.2 ;
          RECT 0.072 0.07 0.09 0.2 ;
          RECT 1.179 0.164 1.197 0.236 ;
          RECT 1.152 0.07 1.197 0.106 ;
          RECT 1.179 0.034 1.197 0.106 ;
          RECT 1.152 0.164 1.197 0.2 ;
          RECT 1.152 0.07 1.17 0.2 ;
          RECT 0.099 0.376 0.117 0.304 ;
          RECT 0.072 0.47 0.117 0.434 ;
          RECT 0.099 0.506 0.117 0.434 ;
          RECT 0.072 0.376 0.117 0.34 ;
          RECT 0.072 0.47 0.09 0.34 ;
          RECT 1.179 0.376 1.197 0.304 ;
          RECT 1.152 0.47 1.197 0.434 ;
          RECT 1.179 0.506 1.197 0.434 ;
          RECT 1.152 0.376 1.197 0.34 ;
          RECT 1.152 0.47 1.17 0.34 ;
          RECT 0.099 0.704 0.117 0.776 ;
          RECT 0.072 0.61 0.117 0.646 ;
          RECT 0.099 0.574 0.117 0.646 ;
          RECT 0.072 0.704 0.117 0.74 ;
          RECT 0.072 0.61 0.09 0.74 ;
          RECT 1.179 0.704 1.197 0.776 ;
          RECT 1.152 0.61 1.197 0.646 ;
          RECT 1.179 0.574 1.197 0.646 ;
          RECT 1.152 0.704 1.197 0.74 ;
          RECT 1.152 0.61 1.17 0.74 ;
          RECT 0.099 0.916 0.117 0.844 ;
          RECT 0.072 1.01 0.117 0.974 ;
          RECT 0.099 1.046 0.117 0.974 ;
          RECT 0.072 0.916 0.117 0.88 ;
          RECT 0.072 1.01 0.09 0.88 ;
          RECT 1.179 0.916 1.197 0.844 ;
          RECT 1.152 1.01 1.197 0.974 ;
          RECT 1.179 1.046 1.197 0.974 ;
          RECT 1.152 0.916 1.197 0.88 ;
          RECT 1.152 1.01 1.17 0.88 ;
          RECT 0.099 1.244 0.117 1.316 ;
          RECT 0.072 1.15 0.117 1.186 ;
          RECT 0.099 1.114 0.117 1.186 ;
          RECT 0.072 1.244 0.117 1.28 ;
          RECT 0.072 1.15 0.09 1.28 ;
          RECT 1.179 1.244 1.197 1.316 ;
          RECT 1.152 1.15 1.197 1.186 ;
          RECT 1.179 1.114 1.197 1.186 ;
          RECT 1.152 1.244 1.197 1.28 ;
          RECT 1.152 1.15 1.17 1.28 ;
          RECT 0.099 1.456 0.117 1.384 ;
          RECT 0.072 1.55 0.117 1.514 ;
          RECT 0.099 1.586 0.117 1.514 ;
          RECT 0.072 1.456 0.117 1.42 ;
          RECT 0.072 1.55 0.09 1.42 ;
          RECT 1.179 1.456 1.197 1.384 ;
          RECT 1.152 1.55 1.197 1.514 ;
          RECT 1.179 1.586 1.197 1.514 ;
          RECT 1.152 1.456 1.197 1.42 ;
          RECT 1.152 1.55 1.17 1.42 ;
          RECT 0.099 1.784 0.117 1.856 ;
          RECT 0.072 1.69 0.117 1.726 ;
          RECT 0.099 1.654 0.117 1.726 ;
          RECT 0.072 1.784 0.117 1.82 ;
          RECT 0.072 1.69 0.09 1.82 ;
          RECT 1.179 1.784 1.197 1.856 ;
          RECT 1.152 1.69 1.197 1.726 ;
          RECT 1.179 1.654 1.197 1.726 ;
          RECT 1.152 1.784 1.197 1.82 ;
          RECT 1.152 1.69 1.17 1.82 ;
          RECT 0.099 1.996 0.117 1.924 ;
          RECT 0.072 2.09 0.117 2.054 ;
          RECT 0.099 2.126 0.117 2.054 ;
          RECT 0.072 1.996 0.117 1.96 ;
          RECT 0.072 2.09 0.09 1.96 ;
          RECT 1.179 1.996 1.197 1.924 ;
          RECT 1.152 2.09 1.197 2.054 ;
          RECT 1.179 2.126 1.197 2.054 ;
          RECT 1.152 1.996 1.197 1.96 ;
          RECT 1.152 2.09 1.17 1.96 ;
        LAYER M2 ;
          RECT 0.072 0.072 1.296 0.09 ;
          RECT 0.072 0.45 1.296 0.468 ;
          RECT 0.072 0.612 1.296 0.63 ;
          RECT 0.072 0.99 1.296 1.008 ;
          RECT 0.072 1.152 1.296 1.17 ;
          RECT 0.072 1.53 1.296 1.548 ;
          RECT 0.072 1.692 1.296 1.71 ;
          RECT 0.072 2.07 1.296 2.088 ;
        LAYER V1 ;
          RECT 0.099 0.072 0.117 0.09 ;
          RECT 1.179 0.072 1.197 0.09 ;
          RECT 0.099 0.45 0.117 0.468 ;
          RECT 1.179 0.45 1.197 0.468 ;
          RECT 0.099 0.612 0.117 0.63 ;
          RECT 1.179 0.612 1.197 0.63 ;
          RECT 0.099 0.99 0.117 1.008 ;
          RECT 1.179 0.99 1.197 1.008 ;
          RECT 0.099 1.152 0.117 1.17 ;
          RECT 1.179 1.152 1.197 1.17 ;
          RECT 0.099 1.53 0.117 1.548 ;
          RECT 1.179 1.53 1.197 1.548 ;
          RECT 0.099 1.692 0.117 1.71 ;
          RECT 1.179 1.692 1.197 1.71 ;
          RECT 0.099 2.07 0.117 2.088 ;
          RECT 1.179 2.07 1.197 2.088 ;
        LAYER M3 ;
          RECT 0.171 0.054 0.189 2.106 ;
        LAYER V2 ;
          RECT 0.171 0.072 0.189 0.09 ;
          RECT 0.171 0.45 0.189 0.468 ;
          RECT 0.171 0.612 0.189 0.63 ;
          RECT 0.171 0.99 0.189 1.008 ;
          RECT 0.171 1.152 0.189 1.17 ;
          RECT 0.171 1.53 0.189 1.548 ;
          RECT 0.171 1.692 0.189 1.71 ;
          RECT 0.171 2.07 0.189 2.088 ;
      END
    END CLK
    PIN D0
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.126 0.29 0.144 ;
          RECT 0.234 0.225 0.271 0.243 ;
          RECT 0.234 0.027 0.271 0.045 ;
          RECT 0.234 0.027 0.252 0.243 ;
      END
    END D0
    PIN QN0
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.225 1.062 0.243 ;
          RECT 1.044 0.027 1.062 0.243 ;
          RECT 1.012 0.027 1.062 0.045 ;
      END
    END QN0
    PIN D1
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 0.126 1.37 0.144 ;
          RECT 1.314 0.225 1.351 0.243 ;
          RECT 1.314 0.027 1.351 0.045 ;
          RECT 1.314 0.027 1.332 0.243 ;
      END
    END D1
    PIN QN1
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 0.225 2.142 0.243 ;
          RECT 2.124 0.027 2.142 0.243 ;
          RECT 2.092 0.027 2.142 0.045 ;
      END
    END QN1
    PIN D2
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.414 0.29 0.396 ;
          RECT 0.234 0.315 0.271 0.297 ;
          RECT 0.234 0.513 0.271 0.495 ;
          RECT 0.234 0.513 0.252 0.297 ;
      END
    END D2
    PIN QN2
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.315 1.062 0.297 ;
          RECT 1.044 0.513 1.062 0.297 ;
          RECT 1.012 0.513 1.062 0.495 ;
      END
    END QN2
    PIN D3
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 0.414 1.37 0.396 ;
          RECT 1.314 0.315 1.351 0.297 ;
          RECT 1.314 0.513 1.351 0.495 ;
          RECT 1.314 0.513 1.332 0.297 ;
      END
    END D3
    PIN QN3
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 0.315 2.142 0.297 ;
          RECT 2.124 0.513 2.142 0.297 ;
          RECT 2.092 0.513 2.142 0.495 ;
      END
    END QN3
    PIN D4
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.666 0.29 0.684 ;
          RECT 0.234 0.765 0.271 0.783 ;
          RECT 0.234 0.567 0.271 0.585 ;
          RECT 0.234 0.567 0.252 0.783 ;
      END
    END D4
    PIN QN4
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.765 1.062 0.783 ;
          RECT 1.044 0.567 1.062 0.783 ;
          RECT 1.012 0.567 1.062 0.585 ;
      END
    END QN4
    PIN D5
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 0.666 1.37 0.684 ;
          RECT 1.314 0.765 1.351 0.783 ;
          RECT 1.314 0.567 1.351 0.585 ;
          RECT 1.314 0.567 1.332 0.783 ;
      END
    END D5
    PIN QN5
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 0.765 2.142 0.783 ;
          RECT 2.124 0.567 2.142 0.783 ;
          RECT 2.092 0.567 2.142 0.585 ;
      END
    END QN5
    PIN D6
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.954 0.29 0.936 ;
          RECT 0.234 0.855 0.271 0.837 ;
          RECT 0.234 1.053 0.271 1.035 ;
          RECT 0.234 1.053 0.252 0.837 ;
      END
    END D6
    PIN QN6
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.855 1.062 0.837 ;
          RECT 1.044 1.053 1.062 0.837 ;
          RECT 1.012 1.053 1.062 1.035 ;
      END
    END QN6
    PIN D7
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 0.954 1.37 0.936 ;
          RECT 1.314 0.855 1.351 0.837 ;
          RECT 1.314 1.053 1.351 1.035 ;
          RECT 1.314 1.053 1.332 0.837 ;
      END
    END D7
    PIN QN7
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 0.855 2.142 0.837 ;
          RECT 2.124 1.053 2.142 0.837 ;
          RECT 2.092 1.053 2.142 1.035 ;
      END
    END QN7
    PIN D8
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.206 0.29 1.224 ;
          RECT 0.234 1.305 0.271 1.323 ;
          RECT 0.234 1.107 0.271 1.125 ;
          RECT 0.234 1.107 0.252 1.323 ;
      END
    END D8
    PIN QN8
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.305 1.062 1.323 ;
          RECT 1.044 1.107 1.062 1.323 ;
          RECT 1.012 1.107 1.062 1.125 ;
      END
    END QN8
    PIN D9
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 1.206 1.37 1.224 ;
          RECT 1.314 1.305 1.351 1.323 ;
          RECT 1.314 1.107 1.351 1.125 ;
          RECT 1.314 1.107 1.332 1.323 ;
      END
    END D9
    PIN QN9
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 1.305 2.142 1.323 ;
          RECT 2.124 1.107 2.142 1.323 ;
          RECT 2.092 1.107 2.142 1.125 ;
      END
    END QN9
    PIN D10
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.494 0.29 1.476 ;
          RECT 0.234 1.395 0.271 1.377 ;
          RECT 0.234 1.593 0.271 1.575 ;
          RECT 0.234 1.593 0.252 1.377 ;
      END
    END D10
    PIN QN10
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.395 1.062 1.377 ;
          RECT 1.044 1.593 1.062 1.377 ;
          RECT 1.012 1.593 1.062 1.575 ;
      END
    END QN10
    PIN D11
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 1.494 1.37 1.476 ;
          RECT 1.314 1.395 1.351 1.377 ;
          RECT 1.314 1.593 1.351 1.575 ;
          RECT 1.314 1.593 1.332 1.377 ;
      END
    END D11
    PIN QN11
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 1.395 2.142 1.377 ;
          RECT 2.124 1.593 2.142 1.377 ;
          RECT 2.092 1.593 2.142 1.575 ;
      END
    END QN11
    PIN D12
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 1.746 0.29 1.764 ;
          RECT 0.234 1.845 0.271 1.863 ;
          RECT 0.234 1.647 0.271 1.665 ;
          RECT 0.234 1.647 0.252 1.863 ;
      END
    END D12
    PIN QN12
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.845 1.062 1.863 ;
          RECT 1.044 1.647 1.062 1.863 ;
          RECT 1.012 1.647 1.062 1.665 ;
      END
    END QN12
    PIN D13
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 1.746 1.37 1.764 ;
          RECT 1.314 1.845 1.351 1.863 ;
          RECT 1.314 1.647 1.351 1.665 ;
          RECT 1.314 1.647 1.332 1.863 ;
      END
    END D13
    PIN QN13
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 1.845 2.142 1.863 ;
          RECT 2.124 1.647 2.142 1.863 ;
          RECT 2.092 1.647 2.142 1.665 ;
      END
    END QN13
    PIN D14
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 2.034 0.29 2.016 ;
          RECT 0.234 1.935 0.271 1.917 ;
          RECT 0.234 2.133 0.271 2.115 ;
          RECT 0.234 2.133 0.252 1.917 ;
      END
    END D14
    PIN QN14
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 1.935 1.062 1.917 ;
          RECT 1.044 2.133 1.062 1.917 ;
          RECT 1.012 2.133 1.062 2.115 ;
      END
    END QN14
    PIN D15
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 1.314 2.034 1.37 2.016 ;
          RECT 1.314 1.935 1.351 1.917 ;
          RECT 1.314 2.133 1.351 2.115 ;
          RECT 1.314 2.133 1.332 1.917 ;
      END
    END D15
    PIN QN15
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 2.092 1.935 2.142 1.917 ;
          RECT 2.124 2.133 2.142 1.917 ;
          RECT 2.092 2.133 2.142 2.115 ;
      END
    END QN15
    OBS
      LAYER M1 ;
        RECT 0.85 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.774 0.027 0.792 0.119 ;
        RECT 0.774 0.027 0.954 0.045 ;
        RECT 0.688 0.224 0.738 0.242 ;
        RECT 0.72 0.027 0.738 0.242 ;
        RECT 0.72 0.153 0.9 0.171 ;
        RECT 0.882 0.117 0.9 0.171 ;
        RECT 0.828 0.117 0.846 0.171 ;
        RECT 0.634 0.027 0.738 0.045 ;
        RECT 0.576 0.225 0.63 0.243 ;
        RECT 0.612 0.081 0.63 0.243 ;
        RECT 0.496 0.081 0.63 0.099 ;
        RECT 0.585 0.045 0.603 0.099 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.45 0.122 0.576 0.14 ;
        RECT 0.418 0.027 0.468 0.045 ;
        RECT 0.315 0.126 0.333 0.203 ;
        RECT 0.315 0.126 0.367 0.144 ;
        RECT 0.148 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.148 0.027 0.198 0.045 ;
        RECT 0.009 0.225 0.068 0.243 ;
        RECT 0.009 0.027 0.027 0.243 ;
        RECT 0.009 0.144 0.047 0.162 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.99 0.09 1.008 0.167 ;
        RECT 0.666 0.101 0.684 0.167 ;
        RECT 0.504 0.165 0.522 0.203 ;
        RECT 0.396 0.106 0.414 0.167 ;
        RECT 0.142 0.106 0.16 0.167 ;
        RECT 1.93 0.225 2.034 0.243 ;
        RECT 2.016 0.027 2.034 0.243 ;
        RECT 1.854 0.027 1.872 0.119 ;
        RECT 1.854 0.027 2.034 0.045 ;
        RECT 1.768 0.224 1.818 0.242 ;
        RECT 1.8 0.027 1.818 0.242 ;
        RECT 1.8 0.153 1.98 0.171 ;
        RECT 1.962 0.117 1.98 0.171 ;
        RECT 1.908 0.117 1.926 0.171 ;
        RECT 1.714 0.027 1.818 0.045 ;
        RECT 1.656 0.225 1.71 0.243 ;
        RECT 1.692 0.081 1.71 0.243 ;
        RECT 1.576 0.081 1.71 0.099 ;
        RECT 1.665 0.045 1.683 0.099 ;
        RECT 1.444 0.225 1.548 0.243 ;
        RECT 1.53 0.027 1.548 0.243 ;
        RECT 1.53 0.122 1.656 0.14 ;
        RECT 1.498 0.027 1.548 0.045 ;
        RECT 1.395 0.126 1.413 0.203 ;
        RECT 1.395 0.126 1.447 0.144 ;
        RECT 1.228 0.225 1.278 0.243 ;
        RECT 1.26 0.027 1.278 0.243 ;
        RECT 1.228 0.027 1.278 0.045 ;
        RECT 1.089 0.225 1.148 0.243 ;
        RECT 1.089 0.027 1.107 0.243 ;
        RECT 1.089 0.144 1.127 0.162 ;
        RECT 1.089 0.027 1.148 0.045 ;
        RECT 2.07 0.09 2.088 0.167 ;
        RECT 1.746 0.101 1.764 0.167 ;
        RECT 1.584 0.165 1.602 0.203 ;
        RECT 1.476 0.106 1.494 0.167 ;
        RECT 1.222 0.106 1.24 0.167 ;
        RECT 0.85 0.315 0.954 0.297 ;
        RECT 0.936 0.513 0.954 0.297 ;
        RECT 0.774 0.513 0.792 0.421 ;
        RECT 0.774 0.513 0.954 0.495 ;
        RECT 0.688 0.316 0.738 0.298 ;
        RECT 0.72 0.513 0.738 0.298 ;
        RECT 0.72 0.387 0.9 0.369 ;
        RECT 0.882 0.423 0.9 0.369 ;
        RECT 0.828 0.423 0.846 0.369 ;
        RECT 0.634 0.513 0.738 0.495 ;
        RECT 0.576 0.315 0.63 0.297 ;
        RECT 0.612 0.459 0.63 0.297 ;
        RECT 0.496 0.459 0.63 0.441 ;
        RECT 0.585 0.495 0.603 0.441 ;
        RECT 0.364 0.315 0.468 0.297 ;
        RECT 0.45 0.513 0.468 0.297 ;
        RECT 0.45 0.418 0.576 0.4 ;
        RECT 0.418 0.513 0.468 0.495 ;
        RECT 0.315 0.414 0.333 0.337 ;
        RECT 0.315 0.414 0.367 0.396 ;
        RECT 0.148 0.315 0.198 0.297 ;
        RECT 0.18 0.513 0.198 0.297 ;
        RECT 0.148 0.513 0.198 0.495 ;
        RECT 0.009 0.315 0.068 0.297 ;
        RECT 0.009 0.513 0.027 0.297 ;
        RECT 0.009 0.396 0.047 0.378 ;
        RECT 0.009 0.513 0.068 0.495 ;
        RECT 0.99 0.45 1.008 0.373 ;
        RECT 0.666 0.439 0.684 0.373 ;
        RECT 0.504 0.375 0.522 0.337 ;
        RECT 0.396 0.434 0.414 0.373 ;
        RECT 0.142 0.434 0.16 0.373 ;
        RECT 1.93 0.315 2.034 0.297 ;
        RECT 2.016 0.513 2.034 0.297 ;
        RECT 1.854 0.513 1.872 0.421 ;
        RECT 1.854 0.513 2.034 0.495 ;
        RECT 1.768 0.316 1.818 0.298 ;
        RECT 1.8 0.513 1.818 0.298 ;
        RECT 1.8 0.387 1.98 0.369 ;
        RECT 1.962 0.423 1.98 0.369 ;
        RECT 1.908 0.423 1.926 0.369 ;
        RECT 1.714 0.513 1.818 0.495 ;
        RECT 1.656 0.315 1.71 0.297 ;
        RECT 1.692 0.459 1.71 0.297 ;
        RECT 1.576 0.459 1.71 0.441 ;
        RECT 1.665 0.495 1.683 0.441 ;
        RECT 1.444 0.315 1.548 0.297 ;
        RECT 1.53 0.513 1.548 0.297 ;
        RECT 1.53 0.418 1.656 0.4 ;
        RECT 1.498 0.513 1.548 0.495 ;
        RECT 1.395 0.414 1.413 0.337 ;
        RECT 1.395 0.414 1.447 0.396 ;
        RECT 1.228 0.315 1.278 0.297 ;
        RECT 1.26 0.513 1.278 0.297 ;
        RECT 1.228 0.513 1.278 0.495 ;
        RECT 1.089 0.315 1.148 0.297 ;
        RECT 1.089 0.513 1.107 0.297 ;
        RECT 1.089 0.396 1.127 0.378 ;
        RECT 1.089 0.513 1.148 0.495 ;
        RECT 2.07 0.45 2.088 0.373 ;
        RECT 1.746 0.439 1.764 0.373 ;
        RECT 1.584 0.375 1.602 0.337 ;
        RECT 1.476 0.434 1.494 0.373 ;
        RECT 1.222 0.434 1.24 0.373 ;
        RECT 0.85 0.765 0.954 0.783 ;
        RECT 0.936 0.567 0.954 0.783 ;
        RECT 0.774 0.567 0.792 0.659 ;
        RECT 0.774 0.567 0.954 0.585 ;
        RECT 0.688 0.764 0.738 0.782 ;
        RECT 0.72 0.567 0.738 0.782 ;
        RECT 0.72 0.693 0.9 0.711 ;
        RECT 0.882 0.657 0.9 0.711 ;
        RECT 0.828 0.657 0.846 0.711 ;
        RECT 0.634 0.567 0.738 0.585 ;
        RECT 0.576 0.765 0.63 0.783 ;
        RECT 0.612 0.621 0.63 0.783 ;
        RECT 0.496 0.621 0.63 0.639 ;
        RECT 0.585 0.585 0.603 0.639 ;
        RECT 0.364 0.765 0.468 0.783 ;
        RECT 0.45 0.567 0.468 0.783 ;
        RECT 0.45 0.662 0.576 0.68 ;
        RECT 0.418 0.567 0.468 0.585 ;
        RECT 0.315 0.666 0.333 0.743 ;
        RECT 0.315 0.666 0.367 0.684 ;
        RECT 0.148 0.765 0.198 0.783 ;
        RECT 0.18 0.567 0.198 0.783 ;
        RECT 0.148 0.567 0.198 0.585 ;
        RECT 0.009 0.765 0.068 0.783 ;
        RECT 0.009 0.567 0.027 0.783 ;
        RECT 0.009 0.684 0.047 0.702 ;
        RECT 0.009 0.567 0.068 0.585 ;
        RECT 0.99 0.63 1.008 0.707 ;
        RECT 0.666 0.641 0.684 0.707 ;
        RECT 0.504 0.705 0.522 0.743 ;
        RECT 0.396 0.646 0.414 0.707 ;
        RECT 0.142 0.646 0.16 0.707 ;
        RECT 1.93 0.765 2.034 0.783 ;
        RECT 2.016 0.567 2.034 0.783 ;
        RECT 1.854 0.567 1.872 0.659 ;
        RECT 1.854 0.567 2.034 0.585 ;
        RECT 1.768 0.764 1.818 0.782 ;
        RECT 1.8 0.567 1.818 0.782 ;
        RECT 1.8 0.693 1.98 0.711 ;
        RECT 1.962 0.657 1.98 0.711 ;
        RECT 1.908 0.657 1.926 0.711 ;
        RECT 1.714 0.567 1.818 0.585 ;
        RECT 1.656 0.765 1.71 0.783 ;
        RECT 1.692 0.621 1.71 0.783 ;
        RECT 1.576 0.621 1.71 0.639 ;
        RECT 1.665 0.585 1.683 0.639 ;
        RECT 1.444 0.765 1.548 0.783 ;
        RECT 1.53 0.567 1.548 0.783 ;
        RECT 1.53 0.662 1.656 0.68 ;
        RECT 1.498 0.567 1.548 0.585 ;
        RECT 1.395 0.666 1.413 0.743 ;
        RECT 1.395 0.666 1.447 0.684 ;
        RECT 1.228 0.765 1.278 0.783 ;
        RECT 1.26 0.567 1.278 0.783 ;
        RECT 1.228 0.567 1.278 0.585 ;
        RECT 1.089 0.765 1.148 0.783 ;
        RECT 1.089 0.567 1.107 0.783 ;
        RECT 1.089 0.684 1.127 0.702 ;
        RECT 1.089 0.567 1.148 0.585 ;
        RECT 2.07 0.63 2.088 0.707 ;
        RECT 1.746 0.641 1.764 0.707 ;
        RECT 1.584 0.705 1.602 0.743 ;
        RECT 1.476 0.646 1.494 0.707 ;
        RECT 1.222 0.646 1.24 0.707 ;
        RECT 0.85 0.855 0.954 0.837 ;
        RECT 0.936 1.053 0.954 0.837 ;
        RECT 0.774 1.053 0.792 0.961 ;
        RECT 0.774 1.053 0.954 1.035 ;
        RECT 0.688 0.856 0.738 0.838 ;
        RECT 0.72 1.053 0.738 0.838 ;
        RECT 0.72 0.927 0.9 0.909 ;
        RECT 0.882 0.963 0.9 0.909 ;
        RECT 0.828 0.963 0.846 0.909 ;
        RECT 0.634 1.053 0.738 1.035 ;
        RECT 0.576 0.855 0.63 0.837 ;
        RECT 0.612 0.999 0.63 0.837 ;
        RECT 0.496 0.999 0.63 0.981 ;
        RECT 0.585 1.035 0.603 0.981 ;
        RECT 0.364 0.855 0.468 0.837 ;
        RECT 0.45 1.053 0.468 0.837 ;
        RECT 0.45 0.958 0.576 0.94 ;
        RECT 0.418 1.053 0.468 1.035 ;
        RECT 0.315 0.954 0.333 0.877 ;
        RECT 0.315 0.954 0.367 0.936 ;
        RECT 0.148 0.855 0.198 0.837 ;
        RECT 0.18 1.053 0.198 0.837 ;
        RECT 0.148 1.053 0.198 1.035 ;
        RECT 0.009 0.855 0.068 0.837 ;
        RECT 0.009 1.053 0.027 0.837 ;
        RECT 0.009 0.936 0.047 0.918 ;
        RECT 0.009 1.053 0.068 1.035 ;
        RECT 0.99 0.99 1.008 0.913 ;
        RECT 0.666 0.979 0.684 0.913 ;
        RECT 0.504 0.915 0.522 0.877 ;
        RECT 0.396 0.974 0.414 0.913 ;
        RECT 0.142 0.974 0.16 0.913 ;
        RECT 1.93 0.855 2.034 0.837 ;
        RECT 2.016 1.053 2.034 0.837 ;
        RECT 1.854 1.053 1.872 0.961 ;
        RECT 1.854 1.053 2.034 1.035 ;
        RECT 1.768 0.856 1.818 0.838 ;
        RECT 1.8 1.053 1.818 0.838 ;
        RECT 1.8 0.927 1.98 0.909 ;
        RECT 1.962 0.963 1.98 0.909 ;
        RECT 1.908 0.963 1.926 0.909 ;
        RECT 1.714 1.053 1.818 1.035 ;
        RECT 1.656 0.855 1.71 0.837 ;
        RECT 1.692 0.999 1.71 0.837 ;
        RECT 1.576 0.999 1.71 0.981 ;
        RECT 1.665 1.035 1.683 0.981 ;
        RECT 1.444 0.855 1.548 0.837 ;
        RECT 1.53 1.053 1.548 0.837 ;
        RECT 1.53 0.958 1.656 0.94 ;
        RECT 1.498 1.053 1.548 1.035 ;
        RECT 1.395 0.954 1.413 0.877 ;
        RECT 1.395 0.954 1.447 0.936 ;
        RECT 1.228 0.855 1.278 0.837 ;
        RECT 1.26 1.053 1.278 0.837 ;
        RECT 1.228 1.053 1.278 1.035 ;
        RECT 1.089 0.855 1.148 0.837 ;
        RECT 1.089 1.053 1.107 0.837 ;
        RECT 1.089 0.936 1.127 0.918 ;
        RECT 1.089 1.053 1.148 1.035 ;
        RECT 2.07 0.99 2.088 0.913 ;
        RECT 1.746 0.979 1.764 0.913 ;
        RECT 1.584 0.915 1.602 0.877 ;
        RECT 1.476 0.974 1.494 0.913 ;
        RECT 1.222 0.974 1.24 0.913 ;
        RECT 0.85 1.305 0.954 1.323 ;
        RECT 0.936 1.107 0.954 1.323 ;
        RECT 0.774 1.107 0.792 1.199 ;
        RECT 0.774 1.107 0.954 1.125 ;
        RECT 0.688 1.304 0.738 1.322 ;
        RECT 0.72 1.107 0.738 1.322 ;
        RECT 0.72 1.233 0.9 1.251 ;
        RECT 0.882 1.197 0.9 1.251 ;
        RECT 0.828 1.197 0.846 1.251 ;
        RECT 0.634 1.107 0.738 1.125 ;
        RECT 0.576 1.305 0.63 1.323 ;
        RECT 0.612 1.161 0.63 1.323 ;
        RECT 0.496 1.161 0.63 1.179 ;
        RECT 0.585 1.125 0.603 1.179 ;
        RECT 0.364 1.305 0.468 1.323 ;
        RECT 0.45 1.107 0.468 1.323 ;
        RECT 0.45 1.202 0.576 1.22 ;
        RECT 0.418 1.107 0.468 1.125 ;
        RECT 0.315 1.206 0.333 1.283 ;
        RECT 0.315 1.206 0.367 1.224 ;
        RECT 0.148 1.305 0.198 1.323 ;
        RECT 0.18 1.107 0.198 1.323 ;
        RECT 0.148 1.107 0.198 1.125 ;
        RECT 0.009 1.305 0.068 1.323 ;
        RECT 0.009 1.107 0.027 1.323 ;
        RECT 0.009 1.224 0.047 1.242 ;
        RECT 0.009 1.107 0.068 1.125 ;
        RECT 0.99 1.17 1.008 1.247 ;
        RECT 0.666 1.181 0.684 1.247 ;
        RECT 0.504 1.245 0.522 1.283 ;
        RECT 0.396 1.186 0.414 1.247 ;
        RECT 0.142 1.186 0.16 1.247 ;
        RECT 1.93 1.305 2.034 1.323 ;
        RECT 2.016 1.107 2.034 1.323 ;
        RECT 1.854 1.107 1.872 1.199 ;
        RECT 1.854 1.107 2.034 1.125 ;
        RECT 1.768 1.304 1.818 1.322 ;
        RECT 1.8 1.107 1.818 1.322 ;
        RECT 1.8 1.233 1.98 1.251 ;
        RECT 1.962 1.197 1.98 1.251 ;
        RECT 1.908 1.197 1.926 1.251 ;
        RECT 1.714 1.107 1.818 1.125 ;
        RECT 1.656 1.305 1.71 1.323 ;
        RECT 1.692 1.161 1.71 1.323 ;
        RECT 1.576 1.161 1.71 1.179 ;
        RECT 1.665 1.125 1.683 1.179 ;
        RECT 1.444 1.305 1.548 1.323 ;
        RECT 1.53 1.107 1.548 1.323 ;
        RECT 1.53 1.202 1.656 1.22 ;
        RECT 1.498 1.107 1.548 1.125 ;
        RECT 1.395 1.206 1.413 1.283 ;
        RECT 1.395 1.206 1.447 1.224 ;
        RECT 1.228 1.305 1.278 1.323 ;
        RECT 1.26 1.107 1.278 1.323 ;
        RECT 1.228 1.107 1.278 1.125 ;
        RECT 1.089 1.305 1.148 1.323 ;
        RECT 1.089 1.107 1.107 1.323 ;
        RECT 1.089 1.224 1.127 1.242 ;
        RECT 1.089 1.107 1.148 1.125 ;
        RECT 2.07 1.17 2.088 1.247 ;
        RECT 1.746 1.181 1.764 1.247 ;
        RECT 1.584 1.245 1.602 1.283 ;
        RECT 1.476 1.186 1.494 1.247 ;
        RECT 1.222 1.186 1.24 1.247 ;
        RECT 0.85 1.395 0.954 1.377 ;
        RECT 0.936 1.593 0.954 1.377 ;
        RECT 0.774 1.593 0.792 1.501 ;
        RECT 0.774 1.593 0.954 1.575 ;
        RECT 0.688 1.396 0.738 1.378 ;
        RECT 0.72 1.593 0.738 1.378 ;
        RECT 0.72 1.467 0.9 1.449 ;
        RECT 0.882 1.503 0.9 1.449 ;
        RECT 0.828 1.503 0.846 1.449 ;
        RECT 0.634 1.593 0.738 1.575 ;
        RECT 0.576 1.395 0.63 1.377 ;
        RECT 0.612 1.539 0.63 1.377 ;
        RECT 0.496 1.539 0.63 1.521 ;
        RECT 0.585 1.575 0.603 1.521 ;
        RECT 0.364 1.395 0.468 1.377 ;
        RECT 0.45 1.593 0.468 1.377 ;
        RECT 0.45 1.498 0.576 1.48 ;
        RECT 0.418 1.593 0.468 1.575 ;
        RECT 0.315 1.494 0.333 1.417 ;
        RECT 0.315 1.494 0.367 1.476 ;
        RECT 0.148 1.395 0.198 1.377 ;
        RECT 0.18 1.593 0.198 1.377 ;
        RECT 0.148 1.593 0.198 1.575 ;
        RECT 0.009 1.395 0.068 1.377 ;
        RECT 0.009 1.593 0.027 1.377 ;
        RECT 0.009 1.476 0.047 1.458 ;
        RECT 0.009 1.593 0.068 1.575 ;
        RECT 0.99 1.53 1.008 1.453 ;
        RECT 0.666 1.519 0.684 1.453 ;
        RECT 0.504 1.455 0.522 1.417 ;
        RECT 0.396 1.514 0.414 1.453 ;
        RECT 0.142 1.514 0.16 1.453 ;
        RECT 1.93 1.395 2.034 1.377 ;
        RECT 2.016 1.593 2.034 1.377 ;
        RECT 1.854 1.593 1.872 1.501 ;
        RECT 1.854 1.593 2.034 1.575 ;
        RECT 1.768 1.396 1.818 1.378 ;
        RECT 1.8 1.593 1.818 1.378 ;
        RECT 1.8 1.467 1.98 1.449 ;
        RECT 1.962 1.503 1.98 1.449 ;
        RECT 1.908 1.503 1.926 1.449 ;
        RECT 1.714 1.593 1.818 1.575 ;
        RECT 1.656 1.395 1.71 1.377 ;
        RECT 1.692 1.539 1.71 1.377 ;
        RECT 1.576 1.539 1.71 1.521 ;
        RECT 1.665 1.575 1.683 1.521 ;
        RECT 1.444 1.395 1.548 1.377 ;
        RECT 1.53 1.593 1.548 1.377 ;
        RECT 1.53 1.498 1.656 1.48 ;
        RECT 1.498 1.593 1.548 1.575 ;
        RECT 1.395 1.494 1.413 1.417 ;
        RECT 1.395 1.494 1.447 1.476 ;
        RECT 1.228 1.395 1.278 1.377 ;
        RECT 1.26 1.593 1.278 1.377 ;
        RECT 1.228 1.593 1.278 1.575 ;
        RECT 1.089 1.395 1.148 1.377 ;
        RECT 1.089 1.593 1.107 1.377 ;
        RECT 1.089 1.476 1.127 1.458 ;
        RECT 1.089 1.593 1.148 1.575 ;
        RECT 2.07 1.53 2.088 1.453 ;
        RECT 1.746 1.519 1.764 1.453 ;
        RECT 1.584 1.455 1.602 1.417 ;
        RECT 1.476 1.514 1.494 1.453 ;
        RECT 1.222 1.514 1.24 1.453 ;
        RECT 0.85 1.845 0.954 1.863 ;
        RECT 0.936 1.647 0.954 1.863 ;
        RECT 0.774 1.647 0.792 1.739 ;
        RECT 0.774 1.647 0.954 1.665 ;
        RECT 0.688 1.844 0.738 1.862 ;
        RECT 0.72 1.647 0.738 1.862 ;
        RECT 0.72 1.773 0.9 1.791 ;
        RECT 0.882 1.737 0.9 1.791 ;
        RECT 0.828 1.737 0.846 1.791 ;
        RECT 0.634 1.647 0.738 1.665 ;
        RECT 0.576 1.845 0.63 1.863 ;
        RECT 0.612 1.701 0.63 1.863 ;
        RECT 0.496 1.701 0.63 1.719 ;
        RECT 0.585 1.665 0.603 1.719 ;
        RECT 0.364 1.845 0.468 1.863 ;
        RECT 0.45 1.647 0.468 1.863 ;
        RECT 0.45 1.742 0.576 1.76 ;
        RECT 0.418 1.647 0.468 1.665 ;
        RECT 0.315 1.746 0.333 1.823 ;
        RECT 0.315 1.746 0.367 1.764 ;
        RECT 0.148 1.845 0.198 1.863 ;
        RECT 0.18 1.647 0.198 1.863 ;
        RECT 0.148 1.647 0.198 1.665 ;
        RECT 0.009 1.845 0.068 1.863 ;
        RECT 0.009 1.647 0.027 1.863 ;
        RECT 0.009 1.764 0.047 1.782 ;
        RECT 0.009 1.647 0.068 1.665 ;
        RECT 0.99 1.71 1.008 1.787 ;
        RECT 0.666 1.721 0.684 1.787 ;
        RECT 0.504 1.785 0.522 1.823 ;
        RECT 0.396 1.726 0.414 1.787 ;
        RECT 0.142 1.726 0.16 1.787 ;
        RECT 1.93 1.845 2.034 1.863 ;
        RECT 2.016 1.647 2.034 1.863 ;
        RECT 1.854 1.647 1.872 1.739 ;
        RECT 1.854 1.647 2.034 1.665 ;
        RECT 1.768 1.844 1.818 1.862 ;
        RECT 1.8 1.647 1.818 1.862 ;
        RECT 1.8 1.773 1.98 1.791 ;
        RECT 1.962 1.737 1.98 1.791 ;
        RECT 1.908 1.737 1.926 1.791 ;
        RECT 1.714 1.647 1.818 1.665 ;
        RECT 1.656 1.845 1.71 1.863 ;
        RECT 1.692 1.701 1.71 1.863 ;
        RECT 1.576 1.701 1.71 1.719 ;
        RECT 1.665 1.665 1.683 1.719 ;
        RECT 1.444 1.845 1.548 1.863 ;
        RECT 1.53 1.647 1.548 1.863 ;
        RECT 1.53 1.742 1.656 1.76 ;
        RECT 1.498 1.647 1.548 1.665 ;
        RECT 1.395 1.746 1.413 1.823 ;
        RECT 1.395 1.746 1.447 1.764 ;
        RECT 1.228 1.845 1.278 1.863 ;
        RECT 1.26 1.647 1.278 1.863 ;
        RECT 1.228 1.647 1.278 1.665 ;
        RECT 1.089 1.845 1.148 1.863 ;
        RECT 1.089 1.647 1.107 1.863 ;
        RECT 1.089 1.764 1.127 1.782 ;
        RECT 1.089 1.647 1.148 1.665 ;
        RECT 2.07 1.71 2.088 1.787 ;
        RECT 1.746 1.721 1.764 1.787 ;
        RECT 1.584 1.785 1.602 1.823 ;
        RECT 1.476 1.726 1.494 1.787 ;
        RECT 1.222 1.726 1.24 1.787 ;
        RECT 0.85 1.935 0.954 1.917 ;
        RECT 0.936 2.133 0.954 1.917 ;
        RECT 0.774 2.133 0.792 2.041 ;
        RECT 0.774 2.133 0.954 2.115 ;
        RECT 0.688 1.936 0.738 1.918 ;
        RECT 0.72 2.133 0.738 1.918 ;
        RECT 0.72 2.007 0.9 1.989 ;
        RECT 0.882 2.043 0.9 1.989 ;
        RECT 0.828 2.043 0.846 1.989 ;
        RECT 0.634 2.133 0.738 2.115 ;
        RECT 0.576 1.935 0.63 1.917 ;
        RECT 0.612 2.079 0.63 1.917 ;
        RECT 0.496 2.079 0.63 2.061 ;
        RECT 0.585 2.115 0.603 2.061 ;
        RECT 0.364 1.935 0.468 1.917 ;
        RECT 0.45 2.133 0.468 1.917 ;
        RECT 0.45 2.038 0.576 2.02 ;
        RECT 0.418 2.133 0.468 2.115 ;
        RECT 0.315 2.034 0.333 1.957 ;
        RECT 0.315 2.034 0.367 2.016 ;
        RECT 0.148 1.935 0.198 1.917 ;
        RECT 0.18 2.133 0.198 1.917 ;
        RECT 0.148 2.133 0.198 2.115 ;
        RECT 0.009 1.935 0.068 1.917 ;
        RECT 0.009 2.133 0.027 1.917 ;
        RECT 0.009 2.016 0.047 1.998 ;
        RECT 0.009 2.133 0.068 2.115 ;
        RECT 0.99 2.07 1.008 1.993 ;
        RECT 0.666 2.059 0.684 1.993 ;
        RECT 0.504 1.995 0.522 1.957 ;
        RECT 0.396 2.054 0.414 1.993 ;
        RECT 0.142 2.054 0.16 1.993 ;
        RECT 1.93 1.935 2.034 1.917 ;
        RECT 2.016 2.133 2.034 1.917 ;
        RECT 1.854 2.133 1.872 2.041 ;
        RECT 1.854 2.133 2.034 2.115 ;
        RECT 1.768 1.936 1.818 1.918 ;
        RECT 1.8 2.133 1.818 1.918 ;
        RECT 1.8 2.007 1.98 1.989 ;
        RECT 1.962 2.043 1.98 1.989 ;
        RECT 1.908 2.043 1.926 1.989 ;
        RECT 1.714 2.133 1.818 2.115 ;
        RECT 1.656 1.935 1.71 1.917 ;
        RECT 1.692 2.079 1.71 1.917 ;
        RECT 1.576 2.079 1.71 2.061 ;
        RECT 1.665 2.115 1.683 2.061 ;
        RECT 1.444 1.935 1.548 1.917 ;
        RECT 1.53 2.133 1.548 1.917 ;
        RECT 1.53 2.038 1.656 2.02 ;
        RECT 1.498 2.133 1.548 2.115 ;
        RECT 1.395 2.034 1.413 1.957 ;
        RECT 1.395 2.034 1.447 2.016 ;
        RECT 1.228 1.935 1.278 1.917 ;
        RECT 1.26 2.133 1.278 1.917 ;
        RECT 1.228 2.133 1.278 2.115 ;
        RECT 1.089 1.935 1.148 1.917 ;
        RECT 1.089 2.133 1.107 1.917 ;
        RECT 1.089 2.016 1.127 1.998 ;
        RECT 1.089 2.133 1.148 2.115 ;
        RECT 2.07 2.07 2.088 1.993 ;
        RECT 1.746 2.059 1.764 1.993 ;
        RECT 1.584 1.995 1.602 1.957 ;
        RECT 1.476 2.054 1.494 1.993 ;
        RECT 1.222 2.054 1.24 1.993 ;
      LAYER M2 ;
        RECT 0.877 0.144 1.013 0.162 ;
        RECT 0.019 0.144 0.689 0.162 ;
        RECT 0.175 0.18 0.527 0.198 ;
        RECT 1.957 0.144 2.093 0.162 ;
        RECT 1.099 0.144 1.769 0.162 ;
        RECT 1.255 0.18 1.607 0.198 ;
        RECT 0.877 0.396 1.013 0.378 ;
        RECT 0.019 0.396 0.689 0.378 ;
        RECT 0.175 0.36 0.527 0.342 ;
        RECT 1.957 0.396 2.093 0.378 ;
        RECT 1.099 0.396 1.769 0.378 ;
        RECT 1.255 0.36 1.607 0.342 ;
        RECT 0.877 0.684 1.013 0.702 ;
        RECT 0.019 0.684 0.689 0.702 ;
        RECT 0.175 0.72 0.527 0.738 ;
        RECT 1.957 0.684 2.093 0.702 ;
        RECT 1.099 0.684 1.769 0.702 ;
        RECT 1.255 0.72 1.607 0.738 ;
        RECT 0.877 0.936 1.013 0.918 ;
        RECT 0.019 0.936 0.689 0.918 ;
        RECT 0.175 0.9 0.527 0.882 ;
        RECT 1.957 0.936 2.093 0.918 ;
        RECT 1.099 0.936 1.769 0.918 ;
        RECT 1.255 0.9 1.607 0.882 ;
        RECT 0.877 1.224 1.013 1.242 ;
        RECT 0.019 1.224 0.689 1.242 ;
        RECT 0.175 1.26 0.527 1.278 ;
        RECT 1.957 1.224 2.093 1.242 ;
        RECT 1.099 1.224 1.769 1.242 ;
        RECT 1.255 1.26 1.607 1.278 ;
        RECT 0.877 1.476 1.013 1.458 ;
        RECT 0.019 1.476 0.689 1.458 ;
        RECT 0.175 1.44 0.527 1.422 ;
        RECT 1.957 1.476 2.093 1.458 ;
        RECT 1.099 1.476 1.769 1.458 ;
        RECT 1.255 1.44 1.607 1.422 ;
        RECT 0.877 1.764 1.013 1.782 ;
        RECT 0.019 1.764 0.689 1.782 ;
        RECT 0.175 1.8 0.527 1.818 ;
        RECT 1.957 1.764 2.093 1.782 ;
        RECT 1.099 1.764 1.769 1.782 ;
        RECT 1.255 1.8 1.607 1.818 ;
        RECT 0.877 2.016 1.013 1.998 ;
        RECT 0.019 2.016 0.689 1.998 ;
        RECT 0.175 1.98 0.527 1.962 ;
        RECT 1.957 2.016 2.093 1.998 ;
        RECT 1.099 2.016 1.769 1.998 ;
        RECT 1.255 1.98 1.607 1.962 ;
      LAYER V1 ;
        RECT 0.99 0.144 1.008 0.162 ;
        RECT 0.882 0.144 0.9 0.162 ;
        RECT 0.666 0.144 0.684 0.162 ;
        RECT 0.504 0.18 0.522 0.198 ;
        RECT 0.396 0.144 0.414 0.162 ;
        RECT 0.315 0.18 0.333 0.198 ;
        RECT 0.18 0.18 0.198 0.198 ;
        RECT 0.142 0.144 0.16 0.162 ;
        RECT 0.024 0.144 0.042 0.162 ;
        RECT 2.07 0.144 2.088 0.162 ;
        RECT 1.962 0.144 1.98 0.162 ;
        RECT 1.746 0.144 1.764 0.162 ;
        RECT 1.584 0.18 1.602 0.198 ;
        RECT 1.476 0.144 1.494 0.162 ;
        RECT 1.395 0.18 1.413 0.198 ;
        RECT 1.26 0.18 1.278 0.198 ;
        RECT 1.222 0.144 1.24 0.162 ;
        RECT 1.104 0.144 1.122 0.162 ;
        RECT 0.99 0.396 1.008 0.378 ;
        RECT 0.882 0.396 0.9 0.378 ;
        RECT 0.666 0.396 0.684 0.378 ;
        RECT 0.504 0.36 0.522 0.342 ;
        RECT 0.396 0.396 0.414 0.378 ;
        RECT 0.315 0.36 0.333 0.342 ;
        RECT 0.18 0.36 0.198 0.342 ;
        RECT 0.142 0.396 0.16 0.378 ;
        RECT 0.024 0.396 0.042 0.378 ;
        RECT 2.07 0.396 2.088 0.378 ;
        RECT 1.962 0.396 1.98 0.378 ;
        RECT 1.746 0.396 1.764 0.378 ;
        RECT 1.584 0.36 1.602 0.342 ;
        RECT 1.476 0.396 1.494 0.378 ;
        RECT 1.395 0.36 1.413 0.342 ;
        RECT 1.26 0.36 1.278 0.342 ;
        RECT 1.222 0.396 1.24 0.378 ;
        RECT 1.104 0.396 1.122 0.378 ;
        RECT 0.99 0.684 1.008 0.702 ;
        RECT 0.882 0.684 0.9 0.702 ;
        RECT 0.666 0.684 0.684 0.702 ;
        RECT 0.504 0.72 0.522 0.738 ;
        RECT 0.396 0.684 0.414 0.702 ;
        RECT 0.315 0.72 0.333 0.738 ;
        RECT 0.18 0.72 0.198 0.738 ;
        RECT 0.142 0.684 0.16 0.702 ;
        RECT 0.024 0.684 0.042 0.702 ;
        RECT 2.07 0.684 2.088 0.702 ;
        RECT 1.962 0.684 1.98 0.702 ;
        RECT 1.746 0.684 1.764 0.702 ;
        RECT 1.584 0.72 1.602 0.738 ;
        RECT 1.476 0.684 1.494 0.702 ;
        RECT 1.395 0.72 1.413 0.738 ;
        RECT 1.26 0.72 1.278 0.738 ;
        RECT 1.222 0.684 1.24 0.702 ;
        RECT 1.104 0.684 1.122 0.702 ;
        RECT 0.99 0.936 1.008 0.918 ;
        RECT 0.882 0.936 0.9 0.918 ;
        RECT 0.666 0.936 0.684 0.918 ;
        RECT 0.504 0.9 0.522 0.882 ;
        RECT 0.396 0.936 0.414 0.918 ;
        RECT 0.315 0.9 0.333 0.882 ;
        RECT 0.18 0.9 0.198 0.882 ;
        RECT 0.142 0.936 0.16 0.918 ;
        RECT 0.024 0.936 0.042 0.918 ;
        RECT 2.07 0.936 2.088 0.918 ;
        RECT 1.962 0.936 1.98 0.918 ;
        RECT 1.746 0.936 1.764 0.918 ;
        RECT 1.584 0.9 1.602 0.882 ;
        RECT 1.476 0.936 1.494 0.918 ;
        RECT 1.395 0.9 1.413 0.882 ;
        RECT 1.26 0.9 1.278 0.882 ;
        RECT 1.222 0.936 1.24 0.918 ;
        RECT 1.104 0.936 1.122 0.918 ;
        RECT 0.99 1.224 1.008 1.242 ;
        RECT 0.882 1.224 0.9 1.242 ;
        RECT 0.666 1.224 0.684 1.242 ;
        RECT 0.504 1.26 0.522 1.278 ;
        RECT 0.396 1.224 0.414 1.242 ;
        RECT 0.315 1.26 0.333 1.278 ;
        RECT 0.18 1.26 0.198 1.278 ;
        RECT 0.142 1.224 0.16 1.242 ;
        RECT 0.024 1.224 0.042 1.242 ;
        RECT 2.07 1.224 2.088 1.242 ;
        RECT 1.962 1.224 1.98 1.242 ;
        RECT 1.746 1.224 1.764 1.242 ;
        RECT 1.584 1.26 1.602 1.278 ;
        RECT 1.476 1.224 1.494 1.242 ;
        RECT 1.395 1.26 1.413 1.278 ;
        RECT 1.26 1.26 1.278 1.278 ;
        RECT 1.222 1.224 1.24 1.242 ;
        RECT 1.104 1.224 1.122 1.242 ;
        RECT 0.99 1.476 1.008 1.458 ;
        RECT 0.882 1.476 0.9 1.458 ;
        RECT 0.666 1.476 0.684 1.458 ;
        RECT 0.504 1.44 0.522 1.422 ;
        RECT 0.396 1.476 0.414 1.458 ;
        RECT 0.315 1.44 0.333 1.422 ;
        RECT 0.18 1.44 0.198 1.422 ;
        RECT 0.142 1.476 0.16 1.458 ;
        RECT 0.024 1.476 0.042 1.458 ;
        RECT 2.07 1.476 2.088 1.458 ;
        RECT 1.962 1.476 1.98 1.458 ;
        RECT 1.746 1.476 1.764 1.458 ;
        RECT 1.584 1.44 1.602 1.422 ;
        RECT 1.476 1.476 1.494 1.458 ;
        RECT 1.395 1.44 1.413 1.422 ;
        RECT 1.26 1.44 1.278 1.422 ;
        RECT 1.222 1.476 1.24 1.458 ;
        RECT 1.104 1.476 1.122 1.458 ;
        RECT 0.99 1.764 1.008 1.782 ;
        RECT 0.882 1.764 0.9 1.782 ;
        RECT 0.666 1.764 0.684 1.782 ;
        RECT 0.504 1.8 0.522 1.818 ;
        RECT 0.396 1.764 0.414 1.782 ;
        RECT 0.315 1.8 0.333 1.818 ;
        RECT 0.18 1.8 0.198 1.818 ;
        RECT 0.142 1.764 0.16 1.782 ;
        RECT 0.024 1.764 0.042 1.782 ;
        RECT 2.07 1.764 2.088 1.782 ;
        RECT 1.962 1.764 1.98 1.782 ;
        RECT 1.746 1.764 1.764 1.782 ;
        RECT 1.584 1.8 1.602 1.818 ;
        RECT 1.476 1.764 1.494 1.782 ;
        RECT 1.395 1.8 1.413 1.818 ;
        RECT 1.26 1.8 1.278 1.818 ;
        RECT 1.222 1.764 1.24 1.782 ;
        RECT 1.104 1.764 1.122 1.782 ;
        RECT 0.99 2.016 1.008 1.998 ;
        RECT 0.882 2.016 0.9 1.998 ;
        RECT 0.666 2.016 0.684 1.998 ;
        RECT 0.504 1.98 0.522 1.962 ;
        RECT 0.396 2.016 0.414 1.998 ;
        RECT 0.315 1.98 0.333 1.962 ;
        RECT 0.18 1.98 0.198 1.962 ;
        RECT 0.142 2.016 0.16 1.998 ;
        RECT 0.024 2.016 0.042 1.998 ;
        RECT 2.07 2.016 2.088 1.998 ;
        RECT 1.962 2.016 1.98 1.998 ;
        RECT 1.746 2.016 1.764 1.998 ;
        RECT 1.584 1.98 1.602 1.962 ;
        RECT 1.476 2.016 1.494 1.998 ;
        RECT 1.395 1.98 1.413 1.962 ;
        RECT 1.26 1.98 1.278 1.962 ;
        RECT 1.222 2.016 1.24 1.998 ;
        RECT 1.104 2.016 1.122 1.998 ;
    END
END DFFHQNV8H2Xx1_ASAP7_75t_L

END LIBRARY
