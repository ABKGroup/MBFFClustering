VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE asap7sc7p5t_R4
  CLASS CORE ;
  SIZE 0.054 BY 1.08 ;
  SYMMETRY Y ;
END asap7sc7p5t_R4

MACRO DFFHQNV4Xx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0.0 0.0 ;
  FOREIGN DFFHQNV4Xx2_ASAP7_75t_L 0.0 0.0 ;
  SIZE 1.134 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_R4 ;
    PIN VDD
      USE POWER ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 0.261 1.134 0.279 ;
          RECT 0.0 0.801 1.134 0.819 ;
      END
    END VDD
    PIN VSS
      USE GROUND ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 -0.009 1.134 0.009 ;
          RECT 0.0 0.549 1.134 0.531 ;
          RECT 0.0 1.089 1.134 1.071 ;
      END
    END VSS
    PIN CLK
      USE CLOCK ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.099 0.164 0.117 0.236 ;
          RECT 0.072 0.07 0.117 0.106 ;
          RECT 0.099 0.034 0.117 0.106 ;
          RECT 0.072 0.164 0.117 0.2 ;
          RECT 0.072 0.07 0.09 0.2 ;
          RECT 0.099 0.376 0.117 0.304 ;
          RECT 0.072 0.47 0.117 0.434 ;
          RECT 0.099 0.506 0.117 0.434 ;
          RECT 0.072 0.376 0.117 0.34 ;
          RECT 0.072 0.47 0.09 0.34 ;
          RECT 0.099 0.704 0.117 0.776 ;
          RECT 0.072 0.61 0.117 0.646 ;
          RECT 0.099 0.574 0.117 0.646 ;
          RECT 0.072 0.704 0.117 0.74 ;
          RECT 0.072 0.61 0.09 0.74 ;
          RECT 0.099 0.916 0.117 0.844 ;
          RECT 0.072 1.01 0.117 0.974 ;
          RECT 0.099 1.046 0.117 0.974 ;
          RECT 0.072 0.916 0.117 0.88 ;
          RECT 0.072 1.01 0.09 0.88 ;
        LAYER M2 ;
          RECT 0.072 0.072 0.216 0.09 ;
          RECT 0.072 0.45 0.216 0.468 ;
          RECT 0.072 0.612 0.216 0.63 ;
          RECT 0.072 0.99 0.216 1.008 ;
        LAYER V1 ;
          RECT 0.099 0.072 0.117 0.09 ;
          RECT 0.099 0.45 0.117 0.468 ;
          RECT 0.099 0.612 0.117 0.63 ;
          RECT 0.099 0.99 0.117 1.008 ;
        LAYER M3 ;
          RECT 0.171 0.054 0.189 1.026 ;
        LAYER V2 ;
          RECT 0.171 0.072 0.189 0.09 ;
          RECT 0.171 0.45 0.189 0.468 ;
          RECT 0.171 0.612 0.189 0.63 ;
          RECT 0.171 0.99 0.189 1.008 ;
      END
    END CLK
    PIN D0
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.126 0.29 0.144 ;
          RECT 0.234 0.225 0.271 0.243 ;
          RECT 0.234 0.027 0.271 0.045 ;
          RECT 0.234 0.027 0.252 0.243 ;
      END
    END D0
    PIN QN0
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.216 1.117 0.234 ;
          RECT 1.099 0.036 1.117 0.234 ;
          RECT 1.012 0.036 1.117 0.054 ;
      END
    END QN0
    PIN D1
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.414 0.29 0.396 ;
          RECT 0.234 0.315 0.271 0.297 ;
          RECT 0.234 0.513 0.271 0.495 ;
          RECT 0.234 0.513 0.252 0.297 ;
      END
    END D1
    PIN QN1
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.324 1.117 0.306 ;
          RECT 1.099 0.504 1.117 0.306 ;
          RECT 1.012 0.504 1.117 0.486 ;
      END
    END QN1
    PIN D2
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.666 0.29 0.684 ;
          RECT 0.234 0.765 0.271 0.783 ;
          RECT 0.234 0.567 0.271 0.585 ;
          RECT 0.234 0.567 0.252 0.783 ;
      END
    END D2
    PIN QN2
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.756 1.117 0.774 ;
          RECT 1.099 0.576 1.117 0.774 ;
          RECT 1.012 0.576 1.117 0.594 ;
      END
    END QN2
    PIN D3
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.954 0.29 0.936 ;
          RECT 0.234 0.855 0.271 0.837 ;
          RECT 0.234 1.053 0.271 1.035 ;
          RECT 0.234 1.053 0.252 0.837 ;
      END
    END D3
    PIN QN3
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.864 1.117 0.846 ;
          RECT 1.099 1.044 1.117 0.846 ;
          RECT 1.012 1.044 1.117 1.026 ;
      END
    END QN3
    OBS
      LAYER M1 ;
        RECT 0.85 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.774 0.027 0.792 0.119 ;
        RECT 0.774 0.027 0.954 0.045 ;
        RECT 0.688 0.224 0.738 0.242 ;
        RECT 0.72 0.027 0.738 0.242 ;
        RECT 0.72 0.153 0.9 0.171 ;
        RECT 0.882 0.117 0.9 0.171 ;
        RECT 0.828 0.117 0.846 0.171 ;
        RECT 0.634 0.027 0.738 0.045 ;
        RECT 0.576 0.225 0.63 0.243 ;
        RECT 0.612 0.081 0.63 0.243 ;
        RECT 0.496 0.081 0.63 0.099 ;
        RECT 0.585 0.045 0.603 0.099 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.45 0.122 0.576 0.14 ;
        RECT 0.418 0.027 0.468 0.045 ;
        RECT 0.315 0.126 0.333 0.203 ;
        RECT 0.315 0.126 0.367 0.144 ;
        RECT 0.148 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.148 0.027 0.198 0.045 ;
        RECT 0.009 0.225 0.068 0.243 ;
        RECT 0.009 0.027 0.027 0.243 ;
        RECT 0.009 0.144 0.047 0.162 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.99 0.09 1.008 0.167 ;
        RECT 0.666 0.101 0.684 0.167 ;
        RECT 0.504 0.165 0.522 0.203 ;
        RECT 0.396 0.106 0.414 0.167 ;
        RECT 0.142 0.106 0.16 0.167 ;
        RECT 0.85 0.315 0.954 0.297 ;
        RECT 0.936 0.513 0.954 0.297 ;
        RECT 0.774 0.513 0.792 0.421 ;
        RECT 0.774 0.513 0.954 0.495 ;
        RECT 0.688 0.316 0.738 0.298 ;
        RECT 0.72 0.513 0.738 0.298 ;
        RECT 0.72 0.387 0.9 0.369 ;
        RECT 0.882 0.423 0.9 0.369 ;
        RECT 0.828 0.423 0.846 0.369 ;
        RECT 0.634 0.513 0.738 0.495 ;
        RECT 0.576 0.315 0.63 0.297 ;
        RECT 0.612 0.459 0.63 0.297 ;
        RECT 0.496 0.459 0.63 0.441 ;
        RECT 0.585 0.495 0.603 0.441 ;
        RECT 0.364 0.315 0.468 0.297 ;
        RECT 0.45 0.513 0.468 0.297 ;
        RECT 0.45 0.418 0.576 0.4 ;
        RECT 0.418 0.513 0.468 0.495 ;
        RECT 0.315 0.414 0.333 0.337 ;
        RECT 0.315 0.414 0.367 0.396 ;
        RECT 0.148 0.315 0.198 0.297 ;
        RECT 0.18 0.513 0.198 0.297 ;
        RECT 0.148 0.513 0.198 0.495 ;
        RECT 0.009 0.315 0.068 0.297 ;
        RECT 0.009 0.513 0.027 0.297 ;
        RECT 0.009 0.396 0.047 0.378 ;
        RECT 0.009 0.513 0.068 0.495 ;
        RECT 0.99 0.45 1.008 0.373 ;
        RECT 0.666 0.439 0.684 0.373 ;
        RECT 0.504 0.375 0.522 0.337 ;
        RECT 0.396 0.434 0.414 0.373 ;
        RECT 0.142 0.434 0.16 0.373 ;
        RECT 0.85 0.765 0.954 0.783 ;
        RECT 0.936 0.567 0.954 0.783 ;
        RECT 0.774 0.567 0.792 0.659 ;
        RECT 0.774 0.567 0.954 0.585 ;
        RECT 0.688 0.764 0.738 0.782 ;
        RECT 0.72 0.567 0.738 0.782 ;
        RECT 0.72 0.693 0.9 0.711 ;
        RECT 0.882 0.657 0.9 0.711 ;
        RECT 0.828 0.657 0.846 0.711 ;
        RECT 0.634 0.567 0.738 0.585 ;
        RECT 0.576 0.765 0.63 0.783 ;
        RECT 0.612 0.621 0.63 0.783 ;
        RECT 0.496 0.621 0.63 0.639 ;
        RECT 0.585 0.585 0.603 0.639 ;
        RECT 0.364 0.765 0.468 0.783 ;
        RECT 0.45 0.567 0.468 0.783 ;
        RECT 0.45 0.662 0.576 0.68 ;
        RECT 0.418 0.567 0.468 0.585 ;
        RECT 0.315 0.666 0.333 0.743 ;
        RECT 0.315 0.666 0.367 0.684 ;
        RECT 0.148 0.765 0.198 0.783 ;
        RECT 0.18 0.567 0.198 0.783 ;
        RECT 0.148 0.567 0.198 0.585 ;
        RECT 0.009 0.765 0.068 0.783 ;
        RECT 0.009 0.567 0.027 0.783 ;
        RECT 0.009 0.684 0.047 0.702 ;
        RECT 0.009 0.567 0.068 0.585 ;
        RECT 0.99 0.63 1.008 0.707 ;
        RECT 0.666 0.641 0.684 0.707 ;
        RECT 0.504 0.705 0.522 0.743 ;
        RECT 0.396 0.646 0.414 0.707 ;
        RECT 0.142 0.646 0.16 0.707 ;
        RECT 0.85 0.855 0.954 0.837 ;
        RECT 0.936 1.053 0.954 0.837 ;
        RECT 0.774 1.053 0.792 0.961 ;
        RECT 0.774 1.053 0.954 1.035 ;
        RECT 0.688 0.856 0.738 0.838 ;
        RECT 0.72 1.053 0.738 0.838 ;
        RECT 0.72 0.927 0.9 0.909 ;
        RECT 0.882 0.963 0.9 0.909 ;
        RECT 0.828 0.963 0.846 0.909 ;
        RECT 0.634 1.053 0.738 1.035 ;
        RECT 0.576 0.855 0.63 0.837 ;
        RECT 0.612 0.999 0.63 0.837 ;
        RECT 0.496 0.999 0.63 0.981 ;
        RECT 0.585 1.035 0.603 0.981 ;
        RECT 0.364 0.855 0.468 0.837 ;
        RECT 0.45 1.053 0.468 0.837 ;
        RECT 0.45 0.958 0.576 0.94 ;
        RECT 0.418 1.053 0.468 1.035 ;
        RECT 0.315 0.954 0.333 0.877 ;
        RECT 0.315 0.954 0.367 0.936 ;
        RECT 0.148 0.855 0.198 0.837 ;
        RECT 0.18 1.053 0.198 0.837 ;
        RECT 0.148 1.053 0.198 1.035 ;
        RECT 0.009 0.855 0.068 0.837 ;
        RECT 0.009 1.053 0.027 0.837 ;
        RECT 0.009 0.936 0.047 0.918 ;
        RECT 0.009 1.053 0.068 1.035 ;
        RECT 0.99 0.99 1.008 0.913 ;
        RECT 0.666 0.979 0.684 0.913 ;
        RECT 0.504 0.915 0.522 0.877 ;
        RECT 0.396 0.974 0.414 0.913 ;
        RECT 0.142 0.974 0.16 0.913 ;
      LAYER M2 ;
        RECT 0.877 0.144 1.013 0.162 ;
        RECT 0.019 0.144 0.689 0.162 ;
        RECT 0.175 0.18 0.527 0.198 ;
        RECT 0.877 0.396 1.013 0.378 ;
        RECT 0.019 0.396 0.689 0.378 ;
        RECT 0.175 0.36 0.527 0.342 ;
        RECT 0.877 0.684 1.013 0.702 ;
        RECT 0.019 0.684 0.689 0.702 ;
        RECT 0.175 0.72 0.527 0.738 ;
        RECT 0.877 0.936 1.013 0.918 ;
        RECT 0.019 0.936 0.689 0.918 ;
        RECT 0.175 0.9 0.527 0.882 ;
      LAYER V1 ;
        RECT 0.99 0.144 1.008 0.162 ;
        RECT 0.882 0.144 0.9 0.162 ;
        RECT 0.666 0.144 0.684 0.162 ;
        RECT 0.504 0.18 0.522 0.198 ;
        RECT 0.396 0.144 0.414 0.162 ;
        RECT 0.315 0.18 0.333 0.198 ;
        RECT 0.18 0.18 0.198 0.198 ;
        RECT 0.142 0.144 0.16 0.162 ;
        RECT 0.024 0.144 0.042 0.162 ;
        RECT 0.99 0.396 1.008 0.378 ;
        RECT 0.882 0.396 0.9 0.378 ;
        RECT 0.666 0.396 0.684 0.378 ;
        RECT 0.504 0.36 0.522 0.342 ;
        RECT 0.396 0.396 0.414 0.378 ;
        RECT 0.315 0.36 0.333 0.342 ;
        RECT 0.18 0.36 0.198 0.342 ;
        RECT 0.142 0.396 0.16 0.378 ;
        RECT 0.024 0.396 0.042 0.378 ;
        RECT 0.99 0.684 1.008 0.702 ;
        RECT 0.882 0.684 0.9 0.702 ;
        RECT 0.666 0.684 0.684 0.702 ;
        RECT 0.504 0.72 0.522 0.738 ;
        RECT 0.396 0.684 0.414 0.702 ;
        RECT 0.315 0.72 0.333 0.738 ;
        RECT 0.18 0.72 0.198 0.738 ;
        RECT 0.142 0.684 0.16 0.702 ;
        RECT 0.024 0.684 0.042 0.702 ;
        RECT 0.99 0.936 1.008 0.918 ;
        RECT 0.882 0.936 0.9 0.918 ;
        RECT 0.666 0.936 0.684 0.918 ;
        RECT 0.504 0.9 0.522 0.882 ;
        RECT 0.396 0.936 0.414 0.918 ;
        RECT 0.315 0.9 0.333 0.882 ;
        RECT 0.18 0.9 0.198 0.882 ;
        RECT 0.142 0.936 0.16 0.918 ;
        RECT 0.024 0.936 0.042 0.918 ;
    END
END DFFHQNV4Xx2_ASAP7_75t_L

END LIBRARY
