VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_256x12
  FOREIGN fakeram7_256x12 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 9.500 BY 11.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.384 0.024 0.408 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.672 0.024 0.696 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.960 0.024 0.984 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.536 0.024 1.560 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.112 0.024 2.136 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.400 0.024 2.424 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.688 0.024 2.712 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.976 0.024 3.000 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.264 0.024 3.288 ;
    END
  END rd_out[11]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.456 0.024 3.480 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.744 0.024 3.768 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.032 0.024 4.056 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.320 0.024 4.344 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.608 0.024 4.632 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.184 0.024 5.208 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.760 0.024 5.784 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 0.024 6.072 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.336 0.024 6.360 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.624 0.024 6.648 ;
    END
  END wd_in[11]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.816 0.024 6.840 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.104 0.024 7.128 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.392 0.024 7.416 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.680 0.024 7.704 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.968 0.024 7.992 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.256 0.024 8.280 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.544 0.024 8.568 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.832 0.024 8.856 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.024 0.024 9.048 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.312 0.024 9.336 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 9.404 0.144 ;
      RECT 0.096 1.584 9.404 1.680 ;
      RECT 0.096 3.120 9.404 3.216 ;
      RECT 0.096 4.656 9.404 4.752 ;
      RECT 0.096 6.192 9.404 6.288 ;
      RECT 0.096 7.728 9.404 7.824 ;
      RECT 0.096 9.264 9.404 9.360 ;
      RECT 0.096 10.800 9.404 10.896 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 9.404 0.912 ;
      RECT 0.096 2.352 9.404 2.448 ;
      RECT 0.096 3.888 9.404 3.984 ;
      RECT 0.096 5.424 9.404 5.520 ;
      RECT 0.096 6.960 9.404 7.056 ;
      RECT 0.096 8.496 9.404 8.592 ;
      RECT 0.096 10.032 9.404 10.128 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 9.500 11.200 ;
    LAYER M2 ;
    RECT 0 0 9.500 11.200 ;
    LAYER M3 ;
    RECT 0 0 9.500 11.200 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 11.200 ;
    RECT 9.404 0 9.500 11.200 ;
    RECT 0.096 0.000 9.404 0.048 ;
    RECT 0.096 0.144 9.404 0.816 ;
    RECT 0.096 0.912 9.404 1.584 ;
    RECT 0.096 1.680 9.404 2.352 ;
    RECT 0.096 2.448 9.404 3.120 ;
    RECT 0.096 3.216 9.404 3.888 ;
    RECT 0.096 3.984 9.404 4.656 ;
    RECT 0.096 4.752 9.404 5.424 ;
    RECT 0.096 5.520 9.404 6.192 ;
    RECT 0.096 6.288 9.404 6.960 ;
    RECT 0.096 7.056 9.404 7.728 ;
    RECT 0.096 7.824 9.404 8.496 ;
    RECT 0.096 8.592 9.404 9.264 ;
    RECT 0.096 9.360 9.404 10.032 ;
    RECT 0.096 10.128 9.404 10.800 ;
    RECT 0.096 10.896 9.404 11.200 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 0.384 ;
    RECT 0 0.408 0.024 0.672 ;
    RECT 0 0.696 0.024 0.960 ;
    RECT 0 0.984 0.024 1.248 ;
    RECT 0 1.272 0.024 1.536 ;
    RECT 0 1.560 0.024 1.824 ;
    RECT 0 1.848 0.024 2.112 ;
    RECT 0 2.136 0.024 2.400 ;
    RECT 0 2.424 0.024 2.688 ;
    RECT 0 2.712 0.024 2.976 ;
    RECT 0 3.000 0.024 3.264 ;
    RECT 0 3.288 0.024 3.456 ;
    RECT 0 3.480 0.024 3.744 ;
    RECT 0 3.768 0.024 4.032 ;
    RECT 0 4.056 0.024 4.320 ;
    RECT 0 4.344 0.024 4.608 ;
    RECT 0 4.632 0.024 4.896 ;
    RECT 0 4.920 0.024 5.184 ;
    RECT 0 5.208 0.024 5.472 ;
    RECT 0 5.496 0.024 5.760 ;
    RECT 0 5.784 0.024 6.048 ;
    RECT 0 6.072 0.024 6.336 ;
    RECT 0 6.360 0.024 6.624 ;
    RECT 0 6.648 0.024 6.816 ;
    RECT 0 6.840 0.024 7.104 ;
    RECT 0 7.128 0.024 7.392 ;
    RECT 0 7.416 0.024 7.680 ;
    RECT 0 7.704 0.024 7.968 ;
    RECT 0 7.992 0.024 8.256 ;
    RECT 0 8.280 0.024 8.544 ;
    RECT 0 8.568 0.024 8.832 ;
    RECT 0 8.856 0.024 9.120 ;
    RECT 0 9.144 0.024 9.408 ;
    RECT 0 9.432 0.024 9.696 ;
    RECT 0 9.720 0.024 9.984 ;
    RECT 0 10.008 0.024 10.176 ;
    RECT 0 10.200 0.024 10.464 ;
    RECT 0 10.488 0.024 10.752 ;
    RECT 0 10.776 0.024 11.040 ;
    RECT 0 11.064 0.024 11.328 ;
    RECT 0 11.352 0.024 11.616 ;
    RECT 0 11.640 0.024 11.904 ;
    RECT 0 11.928 0.024 12.192 ;
    RECT 0 12.216 0.024 12.384 ;
    RECT 0 12.408 0.024 12.672 ;
    RECT 0 12.696 0.024 12.960 ;
    RECT 0 12.984 0.024 11.200 ;
    LAYER OVERLAP ;
    RECT 0 0 9.500 11.200 ;
  END
END fakeram7_256x12

END LIBRARY
