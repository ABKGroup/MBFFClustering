VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_256x32
  FOREIGN fakeram7_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 16.720 BY 16.800 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.288 0.024 0.312 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.480 0.024 0.504 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.672 0.024 0.696 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.864 0.024 0.888 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.056 0.024 1.080 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.632 0.024 1.656 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.016 0.024 2.040 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.208 0.024 2.232 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.400 0.024 2.424 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.592 0.024 2.616 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.784 0.024 2.808 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.976 0.024 3.000 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.360 0.024 3.384 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.552 0.024 3.576 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.744 0.024 3.768 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.936 0.024 3.960 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.320 0.024 4.344 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.512 0.024 4.536 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.704 0.024 4.728 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.088 0.024 5.112 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.280 0.024 5.304 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.664 0.024 5.688 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.856 0.024 5.880 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 0.024 6.072 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.528 0.024 6.552 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.720 0.024 6.744 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.912 0.024 6.936 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.104 0.024 7.128 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.296 0.024 7.320 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.680 0.024 7.704 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.872 0.024 7.896 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.064 0.024 8.088 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.256 0.024 8.280 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.448 0.024 8.472 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.640 0.024 8.664 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.832 0.024 8.856 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.024 0.024 9.048 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.216 0.024 9.240 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.408 0.024 9.432 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.792 0.024 9.816 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.984 0.024 10.008 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.176 0.024 10.200 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.368 0.024 10.392 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.560 0.024 10.584 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.752 0.024 10.776 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.944 0.024 10.968 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.136 0.024 11.160 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.520 0.024 11.544 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.712 0.024 11.736 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.904 0.024 11.928 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.096 0.024 12.120 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.288 0.024 12.312 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.480 0.024 12.504 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.960 0.024 12.984 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.152 0.024 13.176 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.344 0.024 13.368 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.536 0.024 13.560 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.728 0.024 13.752 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.920 0.024 13.944 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.112 0.024 14.136 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.304 0.024 14.328 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.784 0.024 14.808 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.976 0.024 15.000 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.168 0.024 15.192 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 16.624 0.144 ;
      RECT 0.096 1.584 16.624 1.680 ;
      RECT 0.096 3.120 16.624 3.216 ;
      RECT 0.096 4.656 16.624 4.752 ;
      RECT 0.096 6.192 16.624 6.288 ;
      RECT 0.096 7.728 16.624 7.824 ;
      RECT 0.096 9.264 16.624 9.360 ;
      RECT 0.096 10.800 16.624 10.896 ;
      RECT 0.096 12.336 16.624 12.432 ;
      RECT 0.096 13.872 16.624 13.968 ;
      RECT 0.096 15.408 16.624 15.504 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 16.624 0.912 ;
      RECT 0.096 2.352 16.624 2.448 ;
      RECT 0.096 3.888 16.624 3.984 ;
      RECT 0.096 5.424 16.624 5.520 ;
      RECT 0.096 6.960 16.624 7.056 ;
      RECT 0.096 8.496 16.624 8.592 ;
      RECT 0.096 10.032 16.624 10.128 ;
      RECT 0.096 11.568 16.624 11.664 ;
      RECT 0.096 13.104 16.624 13.200 ;
      RECT 0.096 14.640 16.624 14.736 ;
      RECT 0.096 16.176 16.624 16.272 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M2 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M3 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 16.800 ;
    RECT 16.624 0 16.720 16.800 ;
    RECT 0.096 0.000 16.624 0.048 ;
    RECT 0.096 0.144 16.624 0.816 ;
    RECT 0.096 0.912 16.624 1.584 ;
    RECT 0.096 1.680 16.624 2.352 ;
    RECT 0.096 2.448 16.624 3.120 ;
    RECT 0.096 3.216 16.624 3.888 ;
    RECT 0.096 3.984 16.624 4.656 ;
    RECT 0.096 4.752 16.624 5.424 ;
    RECT 0.096 5.520 16.624 6.192 ;
    RECT 0.096 6.288 16.624 6.960 ;
    RECT 0.096 7.056 16.624 7.728 ;
    RECT 0.096 7.824 16.624 8.496 ;
    RECT 0.096 8.592 16.624 9.264 ;
    RECT 0.096 9.360 16.624 10.032 ;
    RECT 0.096 10.128 16.624 10.800 ;
    RECT 0.096 10.896 16.624 11.568 ;
    RECT 0.096 11.664 16.624 12.336 ;
    RECT 0.096 12.432 16.624 13.104 ;
    RECT 0.096 13.200 16.624 13.872 ;
    RECT 0.096 13.968 16.624 14.640 ;
    RECT 0.096 14.736 16.624 15.408 ;
    RECT 0.096 15.504 16.624 16.176 ;
    RECT 0.096 16.272 16.624 16.800 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 0.288 ;
    RECT 0 0.312 0.024 0.480 ;
    RECT 0 0.504 0.024 0.672 ;
    RECT 0 0.696 0.024 0.864 ;
    RECT 0 0.888 0.024 1.056 ;
    RECT 0 1.080 0.024 1.248 ;
    RECT 0 1.272 0.024 1.440 ;
    RECT 0 1.464 0.024 1.632 ;
    RECT 0 1.656 0.024 1.824 ;
    RECT 0 1.848 0.024 2.016 ;
    RECT 0 2.040 0.024 2.208 ;
    RECT 0 2.232 0.024 2.400 ;
    RECT 0 2.424 0.024 2.592 ;
    RECT 0 2.616 0.024 2.784 ;
    RECT 0 2.808 0.024 2.976 ;
    RECT 0 3.000 0.024 3.168 ;
    RECT 0 3.192 0.024 3.360 ;
    RECT 0 3.384 0.024 3.552 ;
    RECT 0 3.576 0.024 3.744 ;
    RECT 0 3.768 0.024 3.936 ;
    RECT 0 3.960 0.024 4.128 ;
    RECT 0 4.152 0.024 4.320 ;
    RECT 0 4.344 0.024 4.512 ;
    RECT 0 4.536 0.024 4.704 ;
    RECT 0 4.728 0.024 4.896 ;
    RECT 0 4.920 0.024 5.088 ;
    RECT 0 5.112 0.024 5.280 ;
    RECT 0 5.304 0.024 5.472 ;
    RECT 0 5.496 0.024 5.664 ;
    RECT 0 5.688 0.024 5.856 ;
    RECT 0 5.880 0.024 6.048 ;
    RECT 0 6.072 0.024 6.528 ;
    RECT 0 6.552 0.024 6.720 ;
    RECT 0 6.744 0.024 6.912 ;
    RECT 0 6.936 0.024 7.104 ;
    RECT 0 7.128 0.024 7.296 ;
    RECT 0 7.320 0.024 7.488 ;
    RECT 0 7.512 0.024 7.680 ;
    RECT 0 7.704 0.024 7.872 ;
    RECT 0 7.896 0.024 8.064 ;
    RECT 0 8.088 0.024 8.256 ;
    RECT 0 8.280 0.024 8.448 ;
    RECT 0 8.472 0.024 8.640 ;
    RECT 0 8.664 0.024 8.832 ;
    RECT 0 8.856 0.024 9.024 ;
    RECT 0 9.048 0.024 9.216 ;
    RECT 0 9.240 0.024 9.408 ;
    RECT 0 9.432 0.024 9.600 ;
    RECT 0 9.624 0.024 9.792 ;
    RECT 0 9.816 0.024 9.984 ;
    RECT 0 10.008 0.024 10.176 ;
    RECT 0 10.200 0.024 10.368 ;
    RECT 0 10.392 0.024 10.560 ;
    RECT 0 10.584 0.024 10.752 ;
    RECT 0 10.776 0.024 10.944 ;
    RECT 0 10.968 0.024 11.136 ;
    RECT 0 11.160 0.024 11.328 ;
    RECT 0 11.352 0.024 11.520 ;
    RECT 0 11.544 0.024 11.712 ;
    RECT 0 11.736 0.024 11.904 ;
    RECT 0 11.928 0.024 12.096 ;
    RECT 0 12.120 0.024 12.288 ;
    RECT 0 12.312 0.024 12.480 ;
    RECT 0 12.504 0.024 12.960 ;
    RECT 0 12.984 0.024 13.152 ;
    RECT 0 13.176 0.024 13.344 ;
    RECT 0 13.368 0.024 13.536 ;
    RECT 0 13.560 0.024 13.728 ;
    RECT 0 13.752 0.024 13.920 ;
    RECT 0 13.944 0.024 14.112 ;
    RECT 0 14.136 0.024 14.304 ;
    RECT 0 14.328 0.024 14.496 ;
    RECT 0 14.520 0.024 14.688 ;
    RECT 0 14.712 0.024 14.880 ;
    RECT 0 14.904 0.024 15.072 ;
    RECT 0 15.096 0.024 15.264 ;
    RECT 0 15.288 0.024 15.456 ;
    RECT 0 15.480 0.024 15.648 ;
    RECT 0 15.672 0.024 15.840 ;
    RECT 0 15.864 0.024 16.032 ;
    RECT 0 16.056 0.024 16.224 ;
    RECT 0 16.248 0.024 16.416 ;
    RECT 0 16.440 0.024 16.608 ;
    RECT 0 16.632 0.024 16.800 ;
    RECT 0 16.824 0.024 16.992 ;
    RECT 0 17.016 0.024 17.184 ;
    RECT 0 17.208 0.024 17.376 ;
    RECT 0 17.400 0.024 17.568 ;
    RECT 0 17.592 0.024 17.760 ;
    RECT 0 17.784 0.024 17.952 ;
    RECT 0 17.976 0.024 18.144 ;
    RECT 0 18.168 0.024 18.336 ;
    RECT 0 18.360 0.024 18.528 ;
    RECT 0 18.552 0.024 18.720 ;
    RECT 0 18.744 0.024 18.912 ;
    RECT 0 18.936 0.024 19.392 ;
    RECT 0 19.416 0.024 19.584 ;
    RECT 0 19.608 0.024 19.776 ;
    RECT 0 19.800 0.024 19.968 ;
    RECT 0 19.992 0.024 20.160 ;
    RECT 0 20.184 0.024 20.352 ;
    RECT 0 20.376 0.024 20.544 ;
    RECT 0 20.568 0.024 20.736 ;
    RECT 0 20.760 0.024 21.216 ;
    RECT 0 21.240 0.024 21.408 ;
    RECT 0 21.432 0.024 21.600 ;
    RECT 0 21.624 0.024 16.800 ;
    LAYER OVERLAP ;
    RECT 0 0 16.720 16.800 ;
  END
END fakeram7_256x32

END LIBRARY
