VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_2048x42
  FOREIGN fakeram7_2048x42 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 21.850 BY 133.000 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.784 0.024 2.808 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.816 0.024 6.840 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.160 0.024 8.184 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.504 0.024 9.528 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.848 0.024 10.872 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.192 0.024 12.216 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.536 0.024 13.560 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.880 0.024 14.904 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.224 0.024 16.248 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.568 0.024 17.592 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.912 0.024 18.936 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.256 0.024 20.280 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.600 0.024 21.624 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.944 0.024 22.968 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.288 0.024 24.312 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.632 0.024 25.656 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.976 0.024 27.000 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.320 0.024 28.344 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.664 0.024 29.688 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.008 0.024 31.032 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.352 0.024 32.376 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.696 0.024 33.720 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.040 0.024 35.064 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.384 0.024 36.408 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.728 0.024 37.752 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.072 0.024 39.096 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.416 0.024 40.440 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.760 0.024 41.784 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.104 0.024 43.128 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.448 0.024 44.472 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.792 0.024 45.816 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.136 0.024 47.160 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.480 0.024 48.504 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.824 0.024 49.848 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.168 0.024 51.192 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.512 0.024 52.536 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.856 0.024 53.880 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.200 0.024 55.224 ;
    END
  END rd_out[41]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.392 0.024 55.416 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.736 0.024 56.760 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.080 0.024 58.104 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.424 0.024 59.448 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.768 0.024 60.792 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.112 0.024 62.136 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.456 0.024 63.480 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 64.800 0.024 64.824 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 66.144 0.024 66.168 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 67.488 0.024 67.512 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 68.832 0.024 68.856 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 70.176 0.024 70.200 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 71.520 0.024 71.544 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 72.864 0.024 72.888 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 74.208 0.024 74.232 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 75.552 0.024 75.576 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 76.896 0.024 76.920 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 78.240 0.024 78.264 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 79.584 0.024 79.608 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 80.928 0.024 80.952 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 82.272 0.024 82.296 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 83.616 0.024 83.640 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 84.960 0.024 84.984 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 86.304 0.024 86.328 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 87.648 0.024 87.672 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 88.992 0.024 89.016 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 90.336 0.024 90.360 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 91.680 0.024 91.704 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 93.024 0.024 93.048 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 94.368 0.024 94.392 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 95.712 0.024 95.736 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 97.056 0.024 97.080 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 98.400 0.024 98.424 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 99.744 0.024 99.768 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 101.088 0.024 101.112 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 102.432 0.024 102.456 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 103.776 0.024 103.800 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 105.120 0.024 105.144 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 106.464 0.024 106.488 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 107.808 0.024 107.832 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 109.152 0.024 109.176 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 110.496 0.024 110.520 ;
    END
  END wd_in[41]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 110.688 0.024 110.712 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 112.032 0.024 112.056 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 113.376 0.024 113.400 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 114.720 0.024 114.744 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 116.064 0.024 116.088 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 117.408 0.024 117.432 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 118.752 0.024 118.776 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 120.096 0.024 120.120 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 121.440 0.024 121.464 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 122.784 0.024 122.808 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 124.128 0.024 124.152 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 124.320 0.024 124.344 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 125.664 0.024 125.688 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 127.008 0.024 127.032 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 21.754 0.144 ;
      RECT 0.096 1.584 21.754 1.680 ;
      RECT 0.096 3.120 21.754 3.216 ;
      RECT 0.096 4.656 21.754 4.752 ;
      RECT 0.096 6.192 21.754 6.288 ;
      RECT 0.096 7.728 21.754 7.824 ;
      RECT 0.096 9.264 21.754 9.360 ;
      RECT 0.096 10.800 21.754 10.896 ;
      RECT 0.096 12.336 21.754 12.432 ;
      RECT 0.096 13.872 21.754 13.968 ;
      RECT 0.096 15.408 21.754 15.504 ;
      RECT 0.096 16.944 21.754 17.040 ;
      RECT 0.096 18.480 21.754 18.576 ;
      RECT 0.096 20.016 21.754 20.112 ;
      RECT 0.096 21.552 21.754 21.648 ;
      RECT 0.096 23.088 21.754 23.184 ;
      RECT 0.096 24.624 21.754 24.720 ;
      RECT 0.096 26.160 21.754 26.256 ;
      RECT 0.096 27.696 21.754 27.792 ;
      RECT 0.096 29.232 21.754 29.328 ;
      RECT 0.096 30.768 21.754 30.864 ;
      RECT 0.096 32.304 21.754 32.400 ;
      RECT 0.096 33.840 21.754 33.936 ;
      RECT 0.096 35.376 21.754 35.472 ;
      RECT 0.096 36.912 21.754 37.008 ;
      RECT 0.096 38.448 21.754 38.544 ;
      RECT 0.096 39.984 21.754 40.080 ;
      RECT 0.096 41.520 21.754 41.616 ;
      RECT 0.096 43.056 21.754 43.152 ;
      RECT 0.096 44.592 21.754 44.688 ;
      RECT 0.096 46.128 21.754 46.224 ;
      RECT 0.096 47.664 21.754 47.760 ;
      RECT 0.096 49.200 21.754 49.296 ;
      RECT 0.096 50.736 21.754 50.832 ;
      RECT 0.096 52.272 21.754 52.368 ;
      RECT 0.096 53.808 21.754 53.904 ;
      RECT 0.096 55.344 21.754 55.440 ;
      RECT 0.096 56.880 21.754 56.976 ;
      RECT 0.096 58.416 21.754 58.512 ;
      RECT 0.096 59.952 21.754 60.048 ;
      RECT 0.096 61.488 21.754 61.584 ;
      RECT 0.096 63.024 21.754 63.120 ;
      RECT 0.096 64.560 21.754 64.656 ;
      RECT 0.096 66.096 21.754 66.192 ;
      RECT 0.096 67.632 21.754 67.728 ;
      RECT 0.096 69.168 21.754 69.264 ;
      RECT 0.096 70.704 21.754 70.800 ;
      RECT 0.096 72.240 21.754 72.336 ;
      RECT 0.096 73.776 21.754 73.872 ;
      RECT 0.096 75.312 21.754 75.408 ;
      RECT 0.096 76.848 21.754 76.944 ;
      RECT 0.096 78.384 21.754 78.480 ;
      RECT 0.096 79.920 21.754 80.016 ;
      RECT 0.096 81.456 21.754 81.552 ;
      RECT 0.096 82.992 21.754 83.088 ;
      RECT 0.096 84.528 21.754 84.624 ;
      RECT 0.096 86.064 21.754 86.160 ;
      RECT 0.096 87.600 21.754 87.696 ;
      RECT 0.096 89.136 21.754 89.232 ;
      RECT 0.096 90.672 21.754 90.768 ;
      RECT 0.096 92.208 21.754 92.304 ;
      RECT 0.096 93.744 21.754 93.840 ;
      RECT 0.096 95.280 21.754 95.376 ;
      RECT 0.096 96.816 21.754 96.912 ;
      RECT 0.096 98.352 21.754 98.448 ;
      RECT 0.096 99.888 21.754 99.984 ;
      RECT 0.096 101.424 21.754 101.520 ;
      RECT 0.096 102.960 21.754 103.056 ;
      RECT 0.096 104.496 21.754 104.592 ;
      RECT 0.096 106.032 21.754 106.128 ;
      RECT 0.096 107.568 21.754 107.664 ;
      RECT 0.096 109.104 21.754 109.200 ;
      RECT 0.096 110.640 21.754 110.736 ;
      RECT 0.096 112.176 21.754 112.272 ;
      RECT 0.096 113.712 21.754 113.808 ;
      RECT 0.096 115.248 21.754 115.344 ;
      RECT 0.096 116.784 21.754 116.880 ;
      RECT 0.096 118.320 21.754 118.416 ;
      RECT 0.096 119.856 21.754 119.952 ;
      RECT 0.096 121.392 21.754 121.488 ;
      RECT 0.096 122.928 21.754 123.024 ;
      RECT 0.096 124.464 21.754 124.560 ;
      RECT 0.096 126.000 21.754 126.096 ;
      RECT 0.096 127.536 21.754 127.632 ;
      RECT 0.096 129.072 21.754 129.168 ;
      RECT 0.096 130.608 21.754 130.704 ;
      RECT 0.096 132.144 21.754 132.240 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 21.754 0.912 ;
      RECT 0.096 2.352 21.754 2.448 ;
      RECT 0.096 3.888 21.754 3.984 ;
      RECT 0.096 5.424 21.754 5.520 ;
      RECT 0.096 6.960 21.754 7.056 ;
      RECT 0.096 8.496 21.754 8.592 ;
      RECT 0.096 10.032 21.754 10.128 ;
      RECT 0.096 11.568 21.754 11.664 ;
      RECT 0.096 13.104 21.754 13.200 ;
      RECT 0.096 14.640 21.754 14.736 ;
      RECT 0.096 16.176 21.754 16.272 ;
      RECT 0.096 17.712 21.754 17.808 ;
      RECT 0.096 19.248 21.754 19.344 ;
      RECT 0.096 20.784 21.754 20.880 ;
      RECT 0.096 22.320 21.754 22.416 ;
      RECT 0.096 23.856 21.754 23.952 ;
      RECT 0.096 25.392 21.754 25.488 ;
      RECT 0.096 26.928 21.754 27.024 ;
      RECT 0.096 28.464 21.754 28.560 ;
      RECT 0.096 30.000 21.754 30.096 ;
      RECT 0.096 31.536 21.754 31.632 ;
      RECT 0.096 33.072 21.754 33.168 ;
      RECT 0.096 34.608 21.754 34.704 ;
      RECT 0.096 36.144 21.754 36.240 ;
      RECT 0.096 37.680 21.754 37.776 ;
      RECT 0.096 39.216 21.754 39.312 ;
      RECT 0.096 40.752 21.754 40.848 ;
      RECT 0.096 42.288 21.754 42.384 ;
      RECT 0.096 43.824 21.754 43.920 ;
      RECT 0.096 45.360 21.754 45.456 ;
      RECT 0.096 46.896 21.754 46.992 ;
      RECT 0.096 48.432 21.754 48.528 ;
      RECT 0.096 49.968 21.754 50.064 ;
      RECT 0.096 51.504 21.754 51.600 ;
      RECT 0.096 53.040 21.754 53.136 ;
      RECT 0.096 54.576 21.754 54.672 ;
      RECT 0.096 56.112 21.754 56.208 ;
      RECT 0.096 57.648 21.754 57.744 ;
      RECT 0.096 59.184 21.754 59.280 ;
      RECT 0.096 60.720 21.754 60.816 ;
      RECT 0.096 62.256 21.754 62.352 ;
      RECT 0.096 63.792 21.754 63.888 ;
      RECT 0.096 65.328 21.754 65.424 ;
      RECT 0.096 66.864 21.754 66.960 ;
      RECT 0.096 68.400 21.754 68.496 ;
      RECT 0.096 69.936 21.754 70.032 ;
      RECT 0.096 71.472 21.754 71.568 ;
      RECT 0.096 73.008 21.754 73.104 ;
      RECT 0.096 74.544 21.754 74.640 ;
      RECT 0.096 76.080 21.754 76.176 ;
      RECT 0.096 77.616 21.754 77.712 ;
      RECT 0.096 79.152 21.754 79.248 ;
      RECT 0.096 80.688 21.754 80.784 ;
      RECT 0.096 82.224 21.754 82.320 ;
      RECT 0.096 83.760 21.754 83.856 ;
      RECT 0.096 85.296 21.754 85.392 ;
      RECT 0.096 86.832 21.754 86.928 ;
      RECT 0.096 88.368 21.754 88.464 ;
      RECT 0.096 89.904 21.754 90.000 ;
      RECT 0.096 91.440 21.754 91.536 ;
      RECT 0.096 92.976 21.754 93.072 ;
      RECT 0.096 94.512 21.754 94.608 ;
      RECT 0.096 96.048 21.754 96.144 ;
      RECT 0.096 97.584 21.754 97.680 ;
      RECT 0.096 99.120 21.754 99.216 ;
      RECT 0.096 100.656 21.754 100.752 ;
      RECT 0.096 102.192 21.754 102.288 ;
      RECT 0.096 103.728 21.754 103.824 ;
      RECT 0.096 105.264 21.754 105.360 ;
      RECT 0.096 106.800 21.754 106.896 ;
      RECT 0.096 108.336 21.754 108.432 ;
      RECT 0.096 109.872 21.754 109.968 ;
      RECT 0.096 111.408 21.754 111.504 ;
      RECT 0.096 112.944 21.754 113.040 ;
      RECT 0.096 114.480 21.754 114.576 ;
      RECT 0.096 116.016 21.754 116.112 ;
      RECT 0.096 117.552 21.754 117.648 ;
      RECT 0.096 119.088 21.754 119.184 ;
      RECT 0.096 120.624 21.754 120.720 ;
      RECT 0.096 122.160 21.754 122.256 ;
      RECT 0.096 123.696 21.754 123.792 ;
      RECT 0.096 125.232 21.754 125.328 ;
      RECT 0.096 126.768 21.754 126.864 ;
      RECT 0.096 128.304 21.754 128.400 ;
      RECT 0.096 129.840 21.754 129.936 ;
      RECT 0.096 131.376 21.754 131.472 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 21.850 133.000 ;
    LAYER M2 ;
    RECT 0 0 21.850 133.000 ;
    LAYER M3 ;
    RECT 0 0 21.850 133.000 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 133.000 ;
    RECT 21.754 0 21.850 133.000 ;
    RECT 0.096 0.000 21.754 0.048 ;
    RECT 0.096 0.144 21.754 0.816 ;
    RECT 0.096 0.912 21.754 1.584 ;
    RECT 0.096 1.680 21.754 2.352 ;
    RECT 0.096 2.448 21.754 3.120 ;
    RECT 0.096 3.216 21.754 3.888 ;
    RECT 0.096 3.984 21.754 4.656 ;
    RECT 0.096 4.752 21.754 5.424 ;
    RECT 0.096 5.520 21.754 6.192 ;
    RECT 0.096 6.288 21.754 6.960 ;
    RECT 0.096 7.056 21.754 7.728 ;
    RECT 0.096 7.824 21.754 8.496 ;
    RECT 0.096 8.592 21.754 9.264 ;
    RECT 0.096 9.360 21.754 10.032 ;
    RECT 0.096 10.128 21.754 10.800 ;
    RECT 0.096 10.896 21.754 11.568 ;
    RECT 0.096 11.664 21.754 12.336 ;
    RECT 0.096 12.432 21.754 13.104 ;
    RECT 0.096 13.200 21.754 13.872 ;
    RECT 0.096 13.968 21.754 14.640 ;
    RECT 0.096 14.736 21.754 15.408 ;
    RECT 0.096 15.504 21.754 16.176 ;
    RECT 0.096 16.272 21.754 16.944 ;
    RECT 0.096 17.040 21.754 17.712 ;
    RECT 0.096 17.808 21.754 18.480 ;
    RECT 0.096 18.576 21.754 19.248 ;
    RECT 0.096 19.344 21.754 20.016 ;
    RECT 0.096 20.112 21.754 20.784 ;
    RECT 0.096 20.880 21.754 21.552 ;
    RECT 0.096 21.648 21.754 22.320 ;
    RECT 0.096 22.416 21.754 23.088 ;
    RECT 0.096 23.184 21.754 23.856 ;
    RECT 0.096 23.952 21.754 24.624 ;
    RECT 0.096 24.720 21.754 25.392 ;
    RECT 0.096 25.488 21.754 26.160 ;
    RECT 0.096 26.256 21.754 26.928 ;
    RECT 0.096 27.024 21.754 27.696 ;
    RECT 0.096 27.792 21.754 28.464 ;
    RECT 0.096 28.560 21.754 29.232 ;
    RECT 0.096 29.328 21.754 30.000 ;
    RECT 0.096 30.096 21.754 30.768 ;
    RECT 0.096 30.864 21.754 31.536 ;
    RECT 0.096 31.632 21.754 32.304 ;
    RECT 0.096 32.400 21.754 33.072 ;
    RECT 0.096 33.168 21.754 33.840 ;
    RECT 0.096 33.936 21.754 34.608 ;
    RECT 0.096 34.704 21.754 35.376 ;
    RECT 0.096 35.472 21.754 36.144 ;
    RECT 0.096 36.240 21.754 36.912 ;
    RECT 0.096 37.008 21.754 37.680 ;
    RECT 0.096 37.776 21.754 38.448 ;
    RECT 0.096 38.544 21.754 39.216 ;
    RECT 0.096 39.312 21.754 39.984 ;
    RECT 0.096 40.080 21.754 40.752 ;
    RECT 0.096 40.848 21.754 41.520 ;
    RECT 0.096 41.616 21.754 42.288 ;
    RECT 0.096 42.384 21.754 43.056 ;
    RECT 0.096 43.152 21.754 43.824 ;
    RECT 0.096 43.920 21.754 44.592 ;
    RECT 0.096 44.688 21.754 45.360 ;
    RECT 0.096 45.456 21.754 46.128 ;
    RECT 0.096 46.224 21.754 46.896 ;
    RECT 0.096 46.992 21.754 47.664 ;
    RECT 0.096 47.760 21.754 48.432 ;
    RECT 0.096 48.528 21.754 49.200 ;
    RECT 0.096 49.296 21.754 49.968 ;
    RECT 0.096 50.064 21.754 50.736 ;
    RECT 0.096 50.832 21.754 51.504 ;
    RECT 0.096 51.600 21.754 52.272 ;
    RECT 0.096 52.368 21.754 53.040 ;
    RECT 0.096 53.136 21.754 53.808 ;
    RECT 0.096 53.904 21.754 54.576 ;
    RECT 0.096 54.672 21.754 55.344 ;
    RECT 0.096 55.440 21.754 56.112 ;
    RECT 0.096 56.208 21.754 56.880 ;
    RECT 0.096 56.976 21.754 57.648 ;
    RECT 0.096 57.744 21.754 58.416 ;
    RECT 0.096 58.512 21.754 59.184 ;
    RECT 0.096 59.280 21.754 59.952 ;
    RECT 0.096 60.048 21.754 60.720 ;
    RECT 0.096 60.816 21.754 61.488 ;
    RECT 0.096 61.584 21.754 62.256 ;
    RECT 0.096 62.352 21.754 63.024 ;
    RECT 0.096 63.120 21.754 63.792 ;
    RECT 0.096 63.888 21.754 64.560 ;
    RECT 0.096 64.656 21.754 65.328 ;
    RECT 0.096 65.424 21.754 66.096 ;
    RECT 0.096 66.192 21.754 66.864 ;
    RECT 0.096 66.960 21.754 67.632 ;
    RECT 0.096 67.728 21.754 68.400 ;
    RECT 0.096 68.496 21.754 69.168 ;
    RECT 0.096 69.264 21.754 69.936 ;
    RECT 0.096 70.032 21.754 70.704 ;
    RECT 0.096 70.800 21.754 71.472 ;
    RECT 0.096 71.568 21.754 72.240 ;
    RECT 0.096 72.336 21.754 73.008 ;
    RECT 0.096 73.104 21.754 73.776 ;
    RECT 0.096 73.872 21.754 74.544 ;
    RECT 0.096 74.640 21.754 75.312 ;
    RECT 0.096 75.408 21.754 76.080 ;
    RECT 0.096 76.176 21.754 76.848 ;
    RECT 0.096 76.944 21.754 77.616 ;
    RECT 0.096 77.712 21.754 78.384 ;
    RECT 0.096 78.480 21.754 79.152 ;
    RECT 0.096 79.248 21.754 79.920 ;
    RECT 0.096 80.016 21.754 80.688 ;
    RECT 0.096 80.784 21.754 81.456 ;
    RECT 0.096 81.552 21.754 82.224 ;
    RECT 0.096 82.320 21.754 82.992 ;
    RECT 0.096 83.088 21.754 83.760 ;
    RECT 0.096 83.856 21.754 84.528 ;
    RECT 0.096 84.624 21.754 85.296 ;
    RECT 0.096 85.392 21.754 86.064 ;
    RECT 0.096 86.160 21.754 86.832 ;
    RECT 0.096 86.928 21.754 87.600 ;
    RECT 0.096 87.696 21.754 88.368 ;
    RECT 0.096 88.464 21.754 89.136 ;
    RECT 0.096 89.232 21.754 89.904 ;
    RECT 0.096 90.000 21.754 90.672 ;
    RECT 0.096 90.768 21.754 91.440 ;
    RECT 0.096 91.536 21.754 92.208 ;
    RECT 0.096 92.304 21.754 92.976 ;
    RECT 0.096 93.072 21.754 93.744 ;
    RECT 0.096 93.840 21.754 94.512 ;
    RECT 0.096 94.608 21.754 95.280 ;
    RECT 0.096 95.376 21.754 96.048 ;
    RECT 0.096 96.144 21.754 96.816 ;
    RECT 0.096 96.912 21.754 97.584 ;
    RECT 0.096 97.680 21.754 98.352 ;
    RECT 0.096 98.448 21.754 99.120 ;
    RECT 0.096 99.216 21.754 99.888 ;
    RECT 0.096 99.984 21.754 100.656 ;
    RECT 0.096 100.752 21.754 101.424 ;
    RECT 0.096 101.520 21.754 102.192 ;
    RECT 0.096 102.288 21.754 102.960 ;
    RECT 0.096 103.056 21.754 103.728 ;
    RECT 0.096 103.824 21.754 104.496 ;
    RECT 0.096 104.592 21.754 105.264 ;
    RECT 0.096 105.360 21.754 106.032 ;
    RECT 0.096 106.128 21.754 106.800 ;
    RECT 0.096 106.896 21.754 107.568 ;
    RECT 0.096 107.664 21.754 108.336 ;
    RECT 0.096 108.432 21.754 109.104 ;
    RECT 0.096 109.200 21.754 109.872 ;
    RECT 0.096 109.968 21.754 110.640 ;
    RECT 0.096 110.736 21.754 111.408 ;
    RECT 0.096 111.504 21.754 112.176 ;
    RECT 0.096 112.272 21.754 112.944 ;
    RECT 0.096 113.040 21.754 113.712 ;
    RECT 0.096 113.808 21.754 114.480 ;
    RECT 0.096 114.576 21.754 115.248 ;
    RECT 0.096 115.344 21.754 116.016 ;
    RECT 0.096 116.112 21.754 116.784 ;
    RECT 0.096 116.880 21.754 117.552 ;
    RECT 0.096 117.648 21.754 118.320 ;
    RECT 0.096 118.416 21.754 119.088 ;
    RECT 0.096 119.184 21.754 119.856 ;
    RECT 0.096 119.952 21.754 120.624 ;
    RECT 0.096 120.720 21.754 121.392 ;
    RECT 0.096 121.488 21.754 122.160 ;
    RECT 0.096 122.256 21.754 122.928 ;
    RECT 0.096 123.024 21.754 123.696 ;
    RECT 0.096 123.792 21.754 124.464 ;
    RECT 0.096 124.560 21.754 125.232 ;
    RECT 0.096 125.328 21.754 126.000 ;
    RECT 0.096 126.096 21.754 126.768 ;
    RECT 0.096 126.864 21.754 127.536 ;
    RECT 0.096 127.632 21.754 128.304 ;
    RECT 0.096 128.400 21.754 129.072 ;
    RECT 0.096 129.168 21.754 129.840 ;
    RECT 0.096 129.936 21.754 130.608 ;
    RECT 0.096 130.704 21.754 131.376 ;
    RECT 0.096 131.472 21.754 132.144 ;
    RECT 0.096 132.240 21.754 133.000 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 1.440 ;
    RECT 0 1.464 0.024 2.784 ;
    RECT 0 2.808 0.024 4.128 ;
    RECT 0 4.152 0.024 5.472 ;
    RECT 0 5.496 0.024 6.816 ;
    RECT 0 6.840 0.024 8.160 ;
    RECT 0 8.184 0.024 9.504 ;
    RECT 0 9.528 0.024 10.848 ;
    RECT 0 10.872 0.024 12.192 ;
    RECT 0 12.216 0.024 13.536 ;
    RECT 0 13.560 0.024 14.880 ;
    RECT 0 14.904 0.024 16.224 ;
    RECT 0 16.248 0.024 17.568 ;
    RECT 0 17.592 0.024 18.912 ;
    RECT 0 18.936 0.024 20.256 ;
    RECT 0 20.280 0.024 21.600 ;
    RECT 0 21.624 0.024 22.944 ;
    RECT 0 22.968 0.024 24.288 ;
    RECT 0 24.312 0.024 25.632 ;
    RECT 0 25.656 0.024 26.976 ;
    RECT 0 27.000 0.024 28.320 ;
    RECT 0 28.344 0.024 29.664 ;
    RECT 0 29.688 0.024 31.008 ;
    RECT 0 31.032 0.024 32.352 ;
    RECT 0 32.376 0.024 33.696 ;
    RECT 0 33.720 0.024 35.040 ;
    RECT 0 35.064 0.024 36.384 ;
    RECT 0 36.408 0.024 37.728 ;
    RECT 0 37.752 0.024 39.072 ;
    RECT 0 39.096 0.024 40.416 ;
    RECT 0 40.440 0.024 41.760 ;
    RECT 0 41.784 0.024 43.104 ;
    RECT 0 43.128 0.024 44.448 ;
    RECT 0 44.472 0.024 45.792 ;
    RECT 0 45.816 0.024 47.136 ;
    RECT 0 47.160 0.024 48.480 ;
    RECT 0 48.504 0.024 49.824 ;
    RECT 0 49.848 0.024 51.168 ;
    RECT 0 51.192 0.024 52.512 ;
    RECT 0 52.536 0.024 53.856 ;
    RECT 0 53.880 0.024 55.200 ;
    RECT 0 55.224 0.024 55.392 ;
    RECT 0 55.416 0.024 56.736 ;
    RECT 0 56.760 0.024 58.080 ;
    RECT 0 58.104 0.024 59.424 ;
    RECT 0 59.448 0.024 60.768 ;
    RECT 0 60.792 0.024 62.112 ;
    RECT 0 62.136 0.024 63.456 ;
    RECT 0 63.480 0.024 64.800 ;
    RECT 0 64.824 0.024 66.144 ;
    RECT 0 66.168 0.024 67.488 ;
    RECT 0 67.512 0.024 68.832 ;
    RECT 0 68.856 0.024 70.176 ;
    RECT 0 70.200 0.024 71.520 ;
    RECT 0 71.544 0.024 72.864 ;
    RECT 0 72.888 0.024 74.208 ;
    RECT 0 74.232 0.024 75.552 ;
    RECT 0 75.576 0.024 76.896 ;
    RECT 0 76.920 0.024 78.240 ;
    RECT 0 78.264 0.024 79.584 ;
    RECT 0 79.608 0.024 80.928 ;
    RECT 0 80.952 0.024 82.272 ;
    RECT 0 82.296 0.024 83.616 ;
    RECT 0 83.640 0.024 84.960 ;
    RECT 0 84.984 0.024 86.304 ;
    RECT 0 86.328 0.024 87.648 ;
    RECT 0 87.672 0.024 88.992 ;
    RECT 0 89.016 0.024 90.336 ;
    RECT 0 90.360 0.024 91.680 ;
    RECT 0 91.704 0.024 93.024 ;
    RECT 0 93.048 0.024 94.368 ;
    RECT 0 94.392 0.024 95.712 ;
    RECT 0 95.736 0.024 97.056 ;
    RECT 0 97.080 0.024 98.400 ;
    RECT 0 98.424 0.024 99.744 ;
    RECT 0 99.768 0.024 101.088 ;
    RECT 0 101.112 0.024 102.432 ;
    RECT 0 102.456 0.024 103.776 ;
    RECT 0 103.800 0.024 105.120 ;
    RECT 0 105.144 0.024 106.464 ;
    RECT 0 106.488 0.024 107.808 ;
    RECT 0 107.832 0.024 109.152 ;
    RECT 0 109.176 0.024 110.496 ;
    RECT 0 110.520 0.024 110.688 ;
    RECT 0 110.712 0.024 112.032 ;
    RECT 0 112.056 0.024 113.376 ;
    RECT 0 113.400 0.024 114.720 ;
    RECT 0 114.744 0.024 116.064 ;
    RECT 0 116.088 0.024 117.408 ;
    RECT 0 117.432 0.024 118.752 ;
    RECT 0 118.776 0.024 120.096 ;
    RECT 0 120.120 0.024 121.440 ;
    RECT 0 121.464 0.024 122.784 ;
    RECT 0 122.808 0.024 124.128 ;
    RECT 0 124.152 0.024 125.472 ;
    RECT 0 125.496 0.024 126.816 ;
    RECT 0 126.840 0.024 128.160 ;
    RECT 0 128.184 0.024 129.504 ;
    RECT 0 129.528 0.024 130.848 ;
    RECT 0 130.872 0.024 132.192 ;
    RECT 0 132.216 0.024 133.536 ;
    RECT 0 133.560 0.024 134.880 ;
    RECT 0 134.904 0.024 136.224 ;
    RECT 0 136.248 0.024 137.568 ;
    RECT 0 137.592 0.024 138.912 ;
    RECT 0 138.936 0.024 140.256 ;
    RECT 0 140.280 0.024 141.600 ;
    RECT 0 141.624 0.024 142.944 ;
    RECT 0 142.968 0.024 144.288 ;
    RECT 0 144.312 0.024 145.632 ;
    RECT 0 145.656 0.024 146.976 ;
    RECT 0 147.000 0.024 148.320 ;
    RECT 0 148.344 0.024 149.664 ;
    RECT 0 149.688 0.024 151.008 ;
    RECT 0 151.032 0.024 152.352 ;
    RECT 0 152.376 0.024 153.696 ;
    RECT 0 153.720 0.024 155.040 ;
    RECT 0 155.064 0.024 156.384 ;
    RECT 0 156.408 0.024 157.728 ;
    RECT 0 157.752 0.024 159.072 ;
    RECT 0 159.096 0.024 160.416 ;
    RECT 0 160.440 0.024 161.760 ;
    RECT 0 161.784 0.024 163.104 ;
    RECT 0 163.128 0.024 164.448 ;
    RECT 0 164.472 0.024 165.792 ;
    RECT 0 165.816 0.024 165.984 ;
    RECT 0 166.008 0.024 167.328 ;
    RECT 0 167.352 0.024 168.672 ;
    RECT 0 168.696 0.024 170.016 ;
    RECT 0 170.040 0.024 171.360 ;
    RECT 0 171.384 0.024 172.704 ;
    RECT 0 172.728 0.024 174.048 ;
    RECT 0 174.072 0.024 175.392 ;
    RECT 0 175.416 0.024 176.736 ;
    RECT 0 176.760 0.024 178.080 ;
    RECT 0 178.104 0.024 179.424 ;
    RECT 0 179.448 0.024 179.616 ;
    RECT 0 179.640 0.024 180.960 ;
    RECT 0 180.984 0.024 182.304 ;
    RECT 0 182.328 0.024 133.000 ;
    LAYER OVERLAP ;
    RECT 0 0 21.850 133.000 ;
  END
END fakeram7_2048x42

END LIBRARY
