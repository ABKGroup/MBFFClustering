VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE asap7sc7p5t_R2
  CLASS CORE ;
  SIZE 0.054 BY 0.54 ;
  SYMMETRY Y ;
END asap7sc7p5t_R2

MACRO DFFHQNV2Xx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0.0 0.0 ;
  FOREIGN DFFHQNV2Xx1_ASAP7_75t_R 0.0 0.0 ;
  SIZE 1.08 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_R2 ;
    PIN VDD
      USE POWER ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 0.261 1.08 0.279 ;
      END
    END VDD
    PIN VSS
      USE GROUND ;
      DIRECTION INOUT ;
      SHAPE ABUTMENT ;
      PORT
        LAYER M1 ;
          RECT 0.0 -0.009 1.08 0.009 ;
          RECT 0.0 0.549 1.08 0.531 ;
      END
    END VSS
    PIN CLK
      USE CLOCK ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.099 0.164 0.117 0.236 ;
          RECT 0.072 0.07 0.117 0.106 ;
          RECT 0.099 0.034 0.117 0.106 ;
          RECT 0.072 0.164 0.117 0.2 ;
          RECT 0.072 0.07 0.09 0.2 ;
          RECT 0.099 0.376 0.117 0.304 ;
          RECT 0.072 0.47 0.117 0.434 ;
          RECT 0.099 0.506 0.117 0.434 ;
          RECT 0.072 0.376 0.117 0.34 ;
          RECT 0.072 0.47 0.09 0.34 ;
        LAYER M2 ;
          RECT 0.072 0.072 0.216 0.09 ;
          RECT 0.072 0.45 0.216 0.468 ;
        LAYER V1 ;
          RECT 0.099 0.072 0.117 0.09 ;
          RECT 0.099 0.45 0.117 0.468 ;
        LAYER M3 ;
          RECT 0.171 0.054 0.189 0.486 ;
        LAYER V2 ;
          RECT 0.171 0.072 0.189 0.09 ;
          RECT 0.171 0.45 0.189 0.468 ;
      END
    END CLK
    PIN D0
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.126 0.29 0.144 ;
          RECT 0.234 0.225 0.271 0.243 ;
          RECT 0.234 0.027 0.271 0.045 ;
          RECT 0.234 0.027 0.252 0.243 ;
      END
    END D0
    PIN QN0
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.225 1.062 0.243 ;
          RECT 1.044 0.027 1.062 0.243 ;
          RECT 1.012 0.027 1.062 0.045 ;
      END
    END QN0
    PIN D1
      USE SIGNAL ;
      DIRECTION INPUT ;
      PORT
        LAYER M1 ;
          RECT 0.234 0.414 0.29 0.396 ;
          RECT 0.234 0.315 0.271 0.297 ;
          RECT 0.234 0.513 0.271 0.495 ;
          RECT 0.234 0.513 0.252 0.297 ;
      END
    END D1
    PIN QN1
      USE SIGNAL ;
      DIRECTION OUTPUT ;
      PORT
        LAYER M1 ;
          RECT 1.012 0.315 1.062 0.297 ;
          RECT 1.044 0.513 1.062 0.297 ;
          RECT 1.012 0.513 1.062 0.495 ;
      END
    END QN1
    OBS
      LAYER M1 ;
        RECT 0.85 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.774 0.027 0.792 0.119 ;
        RECT 0.774 0.027 0.954 0.045 ;
        RECT 0.688 0.224 0.738 0.242 ;
        RECT 0.72 0.027 0.738 0.242 ;
        RECT 0.72 0.153 0.9 0.171 ;
        RECT 0.882 0.117 0.9 0.171 ;
        RECT 0.828 0.117 0.846 0.171 ;
        RECT 0.634 0.027 0.738 0.045 ;
        RECT 0.576 0.225 0.63 0.243 ;
        RECT 0.612 0.081 0.63 0.243 ;
        RECT 0.496 0.081 0.63 0.099 ;
        RECT 0.585 0.045 0.603 0.099 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.45 0.122 0.576 0.14 ;
        RECT 0.418 0.027 0.468 0.045 ;
        RECT 0.315 0.126 0.333 0.203 ;
        RECT 0.315 0.126 0.367 0.144 ;
        RECT 0.148 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.148 0.027 0.198 0.045 ;
        RECT 0.009 0.225 0.068 0.243 ;
        RECT 0.009 0.027 0.027 0.243 ;
        RECT 0.009 0.144 0.047 0.162 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.99 0.09 1.008 0.167 ;
        RECT 0.666 0.101 0.684 0.167 ;
        RECT 0.504 0.165 0.522 0.203 ;
        RECT 0.396 0.106 0.414 0.167 ;
        RECT 0.142 0.106 0.16 0.167 ;
        RECT 0.85 0.315 0.954 0.297 ;
        RECT 0.936 0.513 0.954 0.297 ;
        RECT 0.774 0.513 0.792 0.421 ;
        RECT 0.774 0.513 0.954 0.495 ;
        RECT 0.688 0.316 0.738 0.298 ;
        RECT 0.72 0.513 0.738 0.298 ;
        RECT 0.72 0.387 0.9 0.369 ;
        RECT 0.882 0.423 0.9 0.369 ;
        RECT 0.828 0.423 0.846 0.369 ;
        RECT 0.634 0.513 0.738 0.495 ;
        RECT 0.576 0.315 0.63 0.297 ;
        RECT 0.612 0.459 0.63 0.297 ;
        RECT 0.496 0.459 0.63 0.441 ;
        RECT 0.585 0.495 0.603 0.441 ;
        RECT 0.364 0.315 0.468 0.297 ;
        RECT 0.45 0.513 0.468 0.297 ;
        RECT 0.45 0.418 0.576 0.4 ;
        RECT 0.418 0.513 0.468 0.495 ;
        RECT 0.315 0.414 0.333 0.337 ;
        RECT 0.315 0.414 0.367 0.396 ;
        RECT 0.148 0.315 0.198 0.297 ;
        RECT 0.18 0.513 0.198 0.297 ;
        RECT 0.148 0.513 0.198 0.495 ;
        RECT 0.009 0.315 0.068 0.297 ;
        RECT 0.009 0.513 0.027 0.297 ;
        RECT 0.009 0.396 0.047 0.378 ;
        RECT 0.009 0.513 0.068 0.495 ;
        RECT 0.99 0.45 1.008 0.373 ;
        RECT 0.666 0.439 0.684 0.373 ;
        RECT 0.504 0.375 0.522 0.337 ;
        RECT 0.396 0.434 0.414 0.373 ;
        RECT 0.142 0.434 0.16 0.373 ;
      LAYER M2 ;
        RECT 0.877 0.144 1.013 0.162 ;
        RECT 0.019 0.144 0.689 0.162 ;
        RECT 0.175 0.18 0.527 0.198 ;
        RECT 0.877 0.396 1.013 0.378 ;
        RECT 0.019 0.396 0.689 0.378 ;
        RECT 0.175 0.36 0.527 0.342 ;
      LAYER V1 ;
        RECT 0.99 0.144 1.008 0.162 ;
        RECT 0.882 0.144 0.9 0.162 ;
        RECT 0.666 0.144 0.684 0.162 ;
        RECT 0.504 0.18 0.522 0.198 ;
        RECT 0.396 0.144 0.414 0.162 ;
        RECT 0.315 0.18 0.333 0.198 ;
        RECT 0.18 0.18 0.198 0.198 ;
        RECT 0.142 0.144 0.16 0.162 ;
        RECT 0.024 0.144 0.042 0.162 ;
        RECT 0.99 0.396 1.008 0.378 ;
        RECT 0.882 0.396 0.9 0.378 ;
        RECT 0.666 0.396 0.684 0.378 ;
        RECT 0.504 0.36 0.522 0.342 ;
        RECT 0.396 0.396 0.414 0.378 ;
        RECT 0.315 0.36 0.333 0.342 ;
        RECT 0.18 0.36 0.198 0.342 ;
        RECT 0.142 0.396 0.16 0.378 ;
        RECT 0.024 0.396 0.042 0.378 ;
    END
END DFFHQNV2Xx1_ASAP7_75t_R

END LIBRARY
